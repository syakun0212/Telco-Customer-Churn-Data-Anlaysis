,gender,SeniorCitizen,Partner,Dependents,tenure,PhoneService,MultipleLines,InternetService,OnlineSecurity,OnlineBackup,StreamingTV,StreamingMovies,Contract,PaperlessBilling,PaymentMethod,MonthlyCharges,TotalCharges,Churn,Age,AvgMonthlyGBDownload,AvgMonthlyLongDistanceCharges,CLTV,ChurnValue,City,DeviceProtectionPlan,Gender,InternetType,Latitude,Longitude,Married,MonthlyCharge,NumberofDependents,NumberofReferrals,Offer,Population,PremiumTechSupport,Product/ServiceIssuesReported,ReferredaFriend,StreamingMusic,TenureinMonths,TotalCustomerSvcRequests,TotalExtraDataCharges,TotalLongDistanceCharges,TotalRefunds,TotalRegularCharges,Under30,UnlimitedData,ZipCode
0,0,0,1,0,1,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,29.85,29.85,0,36,10,0.0,3964,0,Los Angeles,0,0,Fiber Optic,33.973616,-118.24902,1,29.85,0,0,Offer E,54492,0,0,0,0,1,2,0.0,0.0,0.0,29.85,0,1,90001
1,1,0,0,0,34,1,0,DSL,1,0,0,0,One year,0,Mailed check,56.95,1889.5,0,46,16,17.09,3441,0,Los Angeles,1,1,Fiber Optic,33.949255,-118.246978,0,56.95,0,0,None,44586,0,0,0,0,34,1,30.23,581.06,0.0,1889.5,0,1,90002
2,1,0,0,0,2,1,0,DSL,1,1,0,0,Month-to-month,1,Mailed check,53.85,108.15,1,37,23,10.47,3239,1,Los Angeles,0,1,Fiber Optic,33.964131,-118.272783,0,56.00400000000001,0,0,None,58198,0,0,0,0,2,4,0.0,20.94,0.0,108.15,0,1,90003
3,1,0,0,0,45,0,No phone service,DSL,1,0,0,0,One year,0,Bank transfer (automatic),42.3,1840.75,0,53,10,0.0,4307,0,Los Angeles,1,1,DSL,34.076259,-118.31071499999999,0,42.3,0,0,None,67852,1,0,0,0,45,4,0.0,0.0,0.0,1840.75,0,1,90004
4,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.7,151.65,1,19,56,9.12,2701,1,Los Angeles,0,0,Cable,34.059281,-118.30742,0,73.528,2,0,None,43019,0,0,0,0,2,0,0.0,18.24,0.0,151.65,1,1,90005
5,0,0,0,0,8,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.65,820.5,1,31,29,12.15,5372,1,Los Angeles,1,0,DSL,34.048013,-118.293953,0,103.636,2,0,None,62784,0,1,0,1,8,2,238.0,97.2,0.0,820.5,0,0,90006
6,1,0,0,1,22,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),89.1,1949.4,0,42,53,29.54,4459,0,Los Angeles,0,1,Fiber Optic,34.027337,-118.28515,0,89.1,3,0,Offer D,45025,0,0,0,0,22,0,0.0,649.88,0.0,1949.4,0,1,90007
7,0,0,0,0,10,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,29.75,301.9,0,42,8,0.0,2013,0,Los Angeles,0,0,Fiber Optic,34.008293,-118.34676599999999,0,29.75,0,0,Offer D,30852,0,0,0,0,10,0,0.0,0.0,0.0,301.9,0,1,90008
8,0,0,1,0,28,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,104.8,3046.05,1,23,52,4.89,5003,1,Los Angeles,1,0,DSL,34.062125,-118.31570900000001,1,108.992,3,0,Offer C,1957,1,1,0,1,28,2,1584.0,136.92,0.0,3046.05,1,0,90010
9,1,0,0,1,62,1,0,DSL,1,1,0,0,One year,0,Bank transfer (automatic),56.15,3487.95,0,48,8,7.96,4529,0,Los Angeles,0,1,Fiber Optic,34.007090000000005,-118.25868100000001,0,56.15,0,0,Offer B,101215,0,0,0,0,62,1,0.0,493.52,0.0,3487.95,0,1,90011
10,1,0,1,1,13,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,49.95,587.45,0,37,22,29.68,5764,0,Los Angeles,0,1,Fiber Optic,34.065875,-118.23872800000001,1,49.95,2,1,Offer D,30596,0,0,1,0,13,3,0.0,385.84,0.0,587.45,0,1,90012
11,1,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),18.95,326.8,0,21,0,32.62,4726,0,Los Angeles,0,1,NA,34.044639000000004,-118.24041299999999,0,18.95,0,0,Offer D,9732,0,0,0,0,16,0,0.0,521.92,0.0,326.8,1,0,90013
12,1,0,1,0,58,1,1,Fiber optic,0,0,1,1,One year,0,Credit card (automatic),100.35,5681.1,0,39,10,5.69,6432,0,Los Angeles,1,1,Fiber Optic,34.043144,-118.251977,1,100.35,0,7,Offer B,3524,0,1,1,1,58,2,0.0,330.0200000000001,0.0,5681.1,0,1,90014
13,1,0,0,0,49,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),103.7,5036.3,1,38,12,44.33,5340,1,Los Angeles,1,1,Cable,34.039224,-118.26629299999999,0,107.848,1,0,None,15140,0,2,0,1,49,2,0.0,2172.17,0.0,5036.3,0,1,90015
14,1,0,0,0,25,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,105.5,2686.05,0,27,48,10.4,5822,0,Los Angeles,1,1,Fiber Optic,34.028331,-118.35433799999998,0,105.5,0,0,None,46984,1,0,0,1,25,0,1289.0,260.0,0.0,2686.05,1,0,90016
15,0,0,1,1,69,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),113.25,7895.15,0,48,3,33.23,5141,0,Los Angeles,1,0,DSL,34.052842,-118.264495,1,113.25,0,7,Offer A,20692,1,0,1,1,69,2,237.0,2292.87,0.0,7895.15,0,0,90017
16,0,0,0,0,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.65,1022.95,0,57,0,22.55,5186,0,Los Angeles,0,0,NA,34.028735,-118.31723600000001,0,20.65,0,0,Offer B,47143,0,0,0,0,52,0,0.0,1172.6,0.0,1022.95,0,0,90018
17,1,0,0,1,71,1,1,Fiber optic,1,0,1,1,Two year,0,Bank transfer (automatic),106.7,7382.25,0,61,7,14.67,4479,0,Los Angeles,1,1,DSL,34.049841,-118.33846000000001,0,106.7,0,0,None,67520,0,0,0,1,71,0,0.0,1041.57,0.0,7382.25,0,1,90019
18,0,0,1,1,10,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),55.2,528.35,1,21,76,9.41,5925,1,San Diego,1,0,Cable,32.898613,-117.202937,1,57.40800000000001,0,6,None,4258,1,0,1,0,10,2,40.15,94.1,0.0,528.35,1,1,92121
19,0,0,0,0,21,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,90.05,1862.9,0,30,73,6.49,5982,0,Los Angeles,1,0,Fiber Optic,34.029043,-118.23950400000001,0,90.05,0,0,Offer D,3012,0,0,0,1,21,0,0.0,136.29,0.0,1862.9,0,1,90021
20,1,1,0,0,1,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,39.65,39.65,1,78,9,0.0,5433,1,Los Angeles,1,1,Fiber Optic,34.02381,-118.156582,0,41.236000000000004,0,0,None,68701,0,0,0,0,1,5,0.0,0.0,0.0,39.65,0,0,90022
21,1,0,1,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.8,202.25,0,45,0,11.04,5279,0,Los Angeles,0,1,NA,34.017697,-118.200577,1,19.8,0,10,Offer D,47487,0,0,1,0,12,0,0.0,132.48,0.0,202.25,0,0,90023
22,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.15,20.15,1,29,0,33.58,4832,1,Los Angeles,0,1,NA,34.066303000000005,-118.435479,0,20.15,0,0,None,44150,0,0,0,0,1,1,0.0,33.58,0.0,20.15,1,0,90024
23,0,0,1,0,58,1,1,DSL,0,1,0,0,Two year,1,Credit card (automatic),59.9,3505.1,0,25,76,48.98,6407,0,Los Angeles,0,0,Fiber Optic,34.046174,-118.44633300000001,1,59.9,0,1,Offer B,41175,1,0,1,0,58,1,2664.0,2840.84,0.0,3505.1,1,0,90025
24,1,0,1,1,49,1,0,DSL,1,1,0,0,Month-to-month,0,Credit card (automatic),59.6,2970.3,0,42,30,5.29,4986,0,Los Angeles,0,1,DSL,34.078990999999995,-118.26380400000001,1,59.6,2,3,Offer B,73686,1,0,1,0,49,2,0.0,259.21,0.0,2970.3,0,1,90026
25,0,0,0,0,30,1,0,DSL,1,1,0,0,Month-to-month,1,Bank transfer (automatic),55.3,1530.6,0,25,27,19.41,2725,0,Los Angeles,0,0,Fiber Optic,34.127194,-118.295647,0,55.3,0,0,None,48727,0,0,0,0,30,2,0.0,582.3,0.0,1530.6,1,1,90027
26,1,0,1,1,47,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.35,4749.15,1,61,18,31.35,5789,1,Los Angeles,0,1,Cable,34.099869,-118.326843,1,103.324,1,1,None,30568,0,1,1,1,47,1,0.0,1473.45,0.0,4749.15,0,1,90028
27,1,0,1,1,1,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,30.2,30.2,1,27,64,0.0,2915,1,Los Angeles,0,1,DSL,34.089953,-118.294824,1,31.408,0,1,None,41713,0,2,1,0,1,3,0.0,0.0,0.0,30.2,1,0,90029
28,1,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),90.25,6369.45,0,36,28,10.92,5974,0,Los Angeles,1,1,Fiber Optic,34.085807,-118.206617,1,90.25,0,9,None,38415,1,0,1,1,72,2,1783.0,786.24,0.0,6369.45,0,0,90031
29,0,0,0,1,17,1,0,DSL,0,0,1,1,Month-to-month,1,Mailed check,64.7,1093.1,1,20,45,40.55,3022,1,Los Angeles,0,0,DSL,34.078821000000005,-118.177576,0,67.28800000000001,0,0,None,46960,0,1,0,1,17,5,0.0,689.3499999999998,0.0,1093.1,1,1,90032
30,0,1,1,0,71,1,1,Fiber optic,1,1,0,0,Two year,1,Credit card (automatic),96.35,6766.95,0,69,12,47.02,5309,0,Los Angeles,1,0,Fiber Optic,34.050197999999995,-118.21094599999999,1,96.35,0,3,None,49431,1,0,1,0,71,0,0.0,3338.42,0.0,6766.95,0,1,90033
31,1,1,1,0,2,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),95.5,181.65,0,79,11,33.1,4449,0,Los Angeles,1,1,Fiber Optic,34.030578000000006,-118.39961299999999,1,95.5,0,10,Offer E,58218,0,0,1,0,2,1,20.0,66.2,0.0,181.65,0,0,90034
32,0,0,1,1,27,1,0,DSL,1,1,0,0,One year,0,Mailed check,66.15,1874.45,0,46,13,40.21,3213,0,Los Angeles,1,0,DSL,34.051809000000006,-118.383843,1,66.15,0,5,None,27799,1,0,1,0,27,0,0.0,1085.67,0.0,1874.45,0,1,90035
33,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.2,20.2,0,35,0,24.48,5526,0,Los Angeles,0,1,NA,34.070291,-118.34919099999999,0,20.2,0,0,Offer E,32901,0,0,0,0,1,0,0.0,24.48,0.0,20.2,0,0,90036
34,1,1,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),45.25,45.25,0,71,12,11.89,3144,0,Los Angeles,0,1,DSL,34.002642,-118.287596,0,45.25,0,0,Offer E,56709,0,0,0,0,1,0,0.0,11.89,0.0,45.25,0,1,90037
35,0,0,1,1,72,1,1,Fiber optic,1,1,1,0,Two year,0,Bank transfer (automatic),99.9,7251.7,0,60,26,23.66,5915,0,Los Angeles,0,0,Fiber Optic,34.088017,-118.327168,1,99.9,0,7,None,32562,1,0,1,0,72,1,1885.0,1703.52,0.0,7251.7,0,0,90038
36,1,0,0,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.7,316.9,1,56,64,12.6,2454,1,Los Angeles,0,1,Cable,34.110845,-118.25959499999999,0,72.488,3,0,None,29310,0,1,0,0,5,1,203.0,63.0,0.0,316.9,0,0,90039
37,0,0,0,0,46,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.8,3548.3,0,19,69,42.44,3395,0,Los Angeles,1,0,Cable,33.994524,-118.149953,0,74.8,0,0,Offer B,9805,0,1,0,0,46,1,2448.0,1952.24,0.0,3548.3,1,0,90040
38,1,0,0,0,34,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.35,3549.25,1,51,31,21.69,2941,1,Los Angeles,1,1,Cable,34.137412,-118.20760700000001,0,110.604,1,0,Offer C,27866,0,0,0,1,34,2,1100.0,737.46,0.0,3549.25,0,0,90041
39,0,0,0,0,11,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),97.85,1105.4,1,48,20,27.57,5674,1,Los Angeles,1,0,Cable,34.11572,-118.19275400000001,0,101.764,2,0,None,64672,0,0,0,1,11,0,221.0,303.27,0.0,1105.4,0,0,90042
40,1,0,1,1,10,1,0,DSL,0,1,0,0,One year,0,Mailed check,49.55,475.7,0,53,7,26.17,2392,0,Los Angeles,0,1,Fiber Optic,33.988543,-118.33408100000001,1,49.55,0,6,Offer D,44764,0,0,1,0,10,2,3.33,261.70000000000005,0.0,475.7,0,1,90043
41,0,0,1,1,70,1,1,DSL,1,1,1,0,Two year,1,Credit card (automatic),69.2,4872.35,0,52,23,29.38,4715,0,Los Angeles,0,0,Fiber Optic,33.952714,-118.292061,1,69.2,0,8,None,87383,0,0,1,0,70,1,112.06,2056.6,0.0,4872.35,0,1,90044
42,0,0,1,1,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.75,418.25,0,28,0,8.74,3646,0,Los Angeles,0,0,NA,33.954017,-118.402447,1,20.75,0,8,Offer D,39334,0,0,1,0,17,0,0.0,148.58,0.0,418.25,1,0,90045
43,0,0,0,0,63,1,1,DSL,1,1,1,0,Two year,1,Credit card (automatic),79.85,4861.45,0,36,17,12.82,4595,0,Los Angeles,1,0,Fiber Optic,34.108455,-118.362081,0,79.85,0,0,Offer B,49839,1,1,0,0,63,2,0.0,807.66,0.0,4861.45,0,1,90046
44,0,0,1,0,13,1,1,DSL,1,1,1,0,Month-to-month,1,Electronic check,76.2,981.45,0,42,29,11.79,2569,0,Los Angeles,0,0,Fiber Optic,33.958149,-118.30844099999999,1,76.2,0,1,Offer D,47107,1,1,1,0,13,2,0.0,153.26999999999995,0.0,981.45,0,1,90047
45,0,0,0,0,49,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.5,3906.7,0,49,24,27.2,6434,0,Los Angeles,0,0,Fiber Optic,34.072945000000004,-118.37267,0,84.5,0,0,Offer B,21739,0,1,0,1,49,1,93.76,1332.8,0.0,3906.7,0,1,90048
46,1,0,0,0,2,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,49.25,97,0,22,71,40.75,3805,0,Los Angeles,0,1,Fiber Optic,34.091829,-118.491244,0,49.25,0,0,None,33523,0,1,0,0,2,1,6.89,81.5,0.0,97.0,1,1,90049
47,0,0,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.65,144.15,1,32,21,5.85,5586,1,Los Angeles,0,0,Cable,33.987945,-118.370442,0,83.876,2,0,None,8115,0,1,0,0,2,2,0.0,11.7,0.0,144.15,0,1,90056
48,1,0,0,0,52,1,1,DSL,1,0,1,1,Two year,1,Credit card (automatic),79.75,4217.8,0,23,73,29.16,4142,0,Los Angeles,0,1,Fiber Optic,34.061918,-118.27793899999999,0,79.75,0,0,Offer B,44004,1,0,0,1,52,2,3079.0,1516.32,0.0,4217.8,1,0,90057
49,0,0,1,1,69,1,1,DSL,1,0,0,0,Two year,1,Credit card (automatic),64.15,4254.1,0,64,17,39.88,5128,0,Los Angeles,1,0,Fiber Optic,34.001616999999996,-118.222274,1,64.15,0,7,None,3642,1,0,1,0,69,2,723.0,2751.7200000000007,0.0,4254.1,0,0,90058
50,0,1,0,0,43,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,90.25,3838.75,0,65,26,12.58,2223,0,Los Angeles,0,0,Fiber Optic,33.927254,-118.249826,0,90.25,0,0,Offer B,38128,0,0,0,0,43,1,998.0,540.94,0.0,3838.75,0,0,90059
51,0,0,0,0,15,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),99.1,1426.4,1,34,22,3.96,2966,1,Los Angeles,0,0,Cable,33.921279999999996,-118.27418600000001,0,103.064,1,0,None,24511,0,1,0,1,15,3,0.0,59.4,0.0,1426.4,0,1,90061
52,0,1,1,0,25,1,1,DSL,1,0,1,0,Month-to-month,1,Credit card (automatic),69.5,1752.65,0,65,2,30.6,3154,0,Los Angeles,0,0,DSL,34.003553000000004,-118.30893300000001,1,69.5,0,9,None,29299,1,0,1,0,25,0,3.51,765.0,0.0,1752.65,0,1,90062
53,0,1,1,0,8,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),80.65,633.3,1,74,19,48.85,5302,1,Los Angeles,0,0,Cable,34.044271,-118.18523700000001,1,83.876,1,1,Offer E,55668,0,0,1,0,8,5,120.0,390.8,0.0,633.3,0,0,90063
54,0,1,1,1,60,1,0,DSL,1,1,0,1,One year,1,Credit card (automatic),74.85,4456.35,0,72,16,48.9,5153,0,Los Angeles,1,0,DSL,34.037251,-118.423573,1,74.85,0,9,Offer B,24505,1,0,1,0,60,0,0.0,2934.0,0.0,4456.35,0,1,90064
55,1,1,0,0,18,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.45,1752.55,1,71,57,11.33,3179,1,Los Angeles,0,1,Fiber Optic,34.108833000000004,-118.22971499999998,0,99.26799999999999,3,0,Offer D,47534,0,0,0,1,18,1,0.0,203.94,45.61,1752.55,0,1,90065
56,0,0,1,1,63,1,1,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),99.65,6311.2,0,44,16,1.43,4572,0,Los Angeles,0,0,Fiber Optic,34.002028,-118.430656,1,99.65,0,2,Offer B,55204,0,0,1,1,63,1,1010.0,90.09,0.0,6311.2,0,0,90066
57,1,1,1,1,66,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,108.45,7076.35,0,77,9,21.79,4582,0,Los Angeles,1,1,Cable,34.057496,-118.413959,1,108.45,0,3,None,2527,1,0,1,0,66,1,637.0,1438.14,0.0,7076.35,0,0,90067
58,0,0,1,1,34,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.95,894.3,0,61,0,25.21,5408,0,Los Angeles,0,0,NA,34.137411,-118.328915,1,24.95,0,10,None,21728,0,0,1,0,34,2,0.0,857.14,0.0,894.3,0,0,90068
59,0,0,0,0,72,1,1,Fiber optic,0,0,1,1,Two year,1,Credit card (automatic),107.5,7853.7,0,40,21,9.47,4708,0,West Hollywood,1,0,DSL,34.093781,-118.38106100000002,0,107.5,0,0,None,20408,1,0,0,1,72,0,1649.0,681.84,0.0,7853.7,0,0,90069
60,0,0,1,0,47,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.5,4707.1,0,34,14,38.15,4488,0,Los Angeles,1,0,Fiber Optic,34.052917,-118.255178,1,100.5,0,3,Offer B,21,0,0,1,1,47,1,0.0,1793.05,0.0,4707.1,0,1,90071
61,1,0,0,0,60,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),89.9,5450.7,0,27,52,42.88,6292,0,Los Angeles,0,1,DSL,34.102084000000005,-118.451629,0,89.9,0,0,Offer B,10470,0,0,0,0,60,3,0.0,2572.8,0.0,5450.7,1,1,90077
62,1,0,1,0,72,0,No phone service,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),42.1,2962,0,36,17,0.0,6091,0,Bell,1,1,DSL,33.970343,-118.17136799999999,1,42.1,0,7,Offer A,105285,0,0,1,0,72,0,50.35,0.0,0.0,2962.0,0,1,90201
63,0,0,1,1,18,1,0,DSL,0,0,0,0,One year,1,Credit card (automatic),54.4,957.1,0,43,7,44.97,4948,0,Beverly Hills,1,0,Fiber Optic,34.099891,-118.41433799999999,1,54.4,0,2,Offer D,21397,1,0,1,0,18,0,67.0,809.46,0.0,957.1,0,0,90210
64,0,0,0,0,9,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,94.4,857.25,1,41,32,27.21,5571,1,Beverly Hills,0,0,Cable,34.063947,-118.38300100000001,0,98.17600000000002,2,0,None,8321,0,0,0,1,9,2,0.0,244.89,0.0,857.25,0,1,90211
65,0,0,0,0,3,1,0,DSL,0,1,1,1,Month-to-month,1,Electronic check,75.3,244.1,0,53,20,38.99,5387,0,Beverly Hills,0,0,Cable,34.062095,-118.401508,0,75.3,0,0,Offer E,11355,1,1,0,1,3,1,0.0,116.97,0.0,244.1,0,1,90212
66,1,0,1,0,47,1,1,Fiber optic,0,1,0,0,One year,1,Electronic check,78.9,3650.35,0,32,30,39.52,3817,0,Compton,0,1,Cable,33.88151,-118.234451,1,78.9,0,8,Offer B,47305,0,0,1,0,47,2,1095.0,1857.44,0.0,3650.35,0,0,90220
67,0,0,0,0,31,1,0,DSL,0,1,1,1,Two year,0,Mailed check,79.2,2497.2,0,61,27,25.57,4984,0,Compton,1,0,Fiber Optic,33.885811,-118.20645900000001,0,79.2,0,0,None,51387,1,0,0,1,31,0,0.0,792.67,0.0,2497.2,0,1,90221
68,0,0,1,1,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.15,930.9,0,37,0,26.95,5849,0,Compton,0,0,NA,33.912246,-118.236773,1,20.15,0,5,Offer B,29825,0,0,1,0,50,0,0.0,1347.5,0.0,930.9,0,0,90222
69,1,0,0,0,10,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,79.85,887.35,0,29,42,48.38,5983,0,Culver City,1,1,Fiber Optic,33.993990999999994,-118.39703999999999,0,79.85,0,0,None,31963,0,0,0,0,10,0,0.0,483.8,0.0,887.35,1,1,90230
70,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,49.05,49.05,0,39,5,25.77,3178,0,Culver City,0,1,Fiber Optic,34.019323,-118.391902,0,49.05,0,0,None,15195,1,1,0,0,1,1,0.0,25.77,0.0,49.05,0,1,90232
71,0,0,1,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,20.4,1090.65,0,24,0,5.65,5482,0,Downey,0,0,NA,33.956228,-118.120993,1,20.4,0,3,Offer B,24908,0,1,1,0,52,1,0.0,293.8,0.0,1090.65,1,0,90240
72,1,1,1,1,64,1,1,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),111.6,7099,0,71,10,16.33,4881,0,Downey,1,1,Fiber Optic,33.940884000000004,-118.128628,1,111.6,0,9,Offer B,40152,1,0,1,0,64,1,710.0,1045.12,0.0,7099.0,0,0,90241
73,1,0,1,1,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.25,1424.6,0,40,0,48.73,4444,0,Downey,0,1,NA,33.921793,-118.140588,1,24.25,0,4,Offer B,42459,0,1,1,0,62,1,0.0,3021.26,0.0,1424.6,0,0,90242
74,0,0,0,1,3,1,0,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),64.5,177.4,0,51,56,39.55,5613,0,El Segundo,0,0,Fiber Optic,33.917145,-118.401554,0,64.5,3,0,Offer E,16041,1,0,0,1,3,0,0.0,118.65,0.0,177.4,0,1,90245
75,0,1,0,0,56,1,1,Fiber optic,1,1,1,1,One year,0,Electronic check,110.5,6139.5,0,73,29,47.13,4463,0,Gardena,1,0,Cable,33.890853,-118.29796699999999,0,110.5,0,0,None,47758,0,0,0,0,56,2,0.0,2639.28,0.0,6139.5,0,1,90247
76,0,0,0,0,46,1,0,DSL,0,0,0,1,One year,0,Credit card (automatic),55.65,2688.85,0,50,7,2.03,2867,0,Gardena,0,0,Fiber Optic,33.876482,-118.284077,0,55.65,0,0,Offer B,9960,0,0,0,1,46,0,0.0,93.38,0.0,2688.85,0,1,90248
77,0,0,1,1,8,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,54.65,482.25,0,62,18,38.78,5614,0,Gardena,0,0,Fiber Optic,33.90139,-118.315697,1,54.65,1,1,Offer E,26442,0,0,1,0,8,0,0.0,310.24,0.0,482.25,0,1,90249
78,1,1,0,0,30,1,0,DSL,1,1,1,1,Month-to-month,1,Electronic check,74.75,2111.3,0,80,5,38.61,3033,0,Hawthorne,0,1,DSL,33.914775,-118.348083,0,74.75,0,0,None,93315,0,0,0,0,30,1,106.0,1158.3,0.0,2111.3,0,0,90250
79,0,0,1,1,45,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),25.9,1216.6,0,48,0,22.49,5741,0,Hermosa Beach,0,0,NA,33.865320000000004,-118.396336,1,25.9,0,4,Offer B,18693,0,2,1,0,45,3,0.0,1012.05,0.0,1216.6,0,0,90254
80,0,0,0,1,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.35,79.35,1,32,63,13.13,2483,1,Huntington Park,0,0,Cable,33.97803,-118.217141,0,82.524,3,0,None,78114,0,1,0,0,1,3,0.0,13.13,0.0,79.35,0,0,90255
81,0,0,1,1,11,0,No phone service,DSL,1,0,1,1,Month-to-month,0,Electronic check,50.55,565.35,0,23,41,0.0,3443,0,Lawndale,0,0,Cable,33.88856,-118.35181299999999,1,50.55,1,1,None,33300,0,2,1,1,11,3,23.18,0.0,0.0,565.35,1,1,90260
82,0,0,1,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.15,496.9,1,34,58,8.69,3457,1,Lynwood,1,0,Cable,33.923573,-118.20066899999999,1,78.156,5,1,None,69850,0,0,1,0,7,0,288.0,60.83,0.0,496.9,0,0,90262
83,0,0,0,0,42,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),103.8,4327.5,0,38,28,40.15,4005,0,Malibu,1,0,DSL,34.037037,-118.705803,0,103.8,0,0,Offer B,11,1,0,0,1,42,1,0.0,1686.3,0.0,4327.5,0,1,90263
84,0,0,1,0,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.15,973.35,0,31,0,2.82,5422,0,Malibu,0,0,NA,34.074571999999996,-118.831181,1,20.15,0,10,None,19630,0,0,1,0,49,0,0.0,138.17999999999998,0.0,973.35,0,0,90265
85,1,0,0,0,9,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),99.3,918.75,0,30,69,4.81,3540,0,Manhattan Beach,0,1,DSL,33.889632,-118.39737,0,99.3,0,0,Offer E,33758,0,0,0,1,9,2,634.0,43.29,0.0,918.75,0,0,90266
86,0,0,1,0,35,1,0,DSL,1,0,1,0,One year,1,Bank transfer (automatic),62.15,2215.45,0,51,30,24.53,5255,0,Maywood,0,0,DSL,33.988572,-118.18656499999999,1,62.15,0,1,Offer C,28094,0,0,1,0,35,1,665.0,858.5500000000002,0.0,2215.45,0,0,90270
87,0,0,1,1,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.65,1057,0,24,0,37.96,4124,0,Pacific Palisades,0,0,NA,34.079449,-118.54830600000001,1,20.65,0,10,None,22548,0,0,1,0,48,0,0.0,1822.08,0.0,1057.0,1,0,90272
88,0,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.95,927.1,0,56,0,30.47,5480,0,Palos Verdes Peninsula,0,0,NA,33.788208000000004,-118.404955,1,19.95,0,1,None,24979,0,0,1,0,46,0,0.0,1401.62,0.0,927.1,0,0,90274
89,1,0,1,0,29,0,No phone service,DSL,0,0,1,0,Month-to-month,0,Mailed check,33.75,1009.25,0,47,22,0.0,3664,0,Rancho Palos Verdes,0,1,DSL,33.753146,-118.36745900000001,1,33.75,0,4,Offer C,41263,0,0,1,0,29,0,0.0,0.0,0.0,1009.25,0,1,90275
90,1,0,1,1,30,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),82.05,2570.2,0,32,21,6.19,5036,0,Redondo Beach,1,1,Cable,33.830453000000006,-118.384565,1,82.05,3,5,Offer C,34191,0,0,1,0,30,0,540.0,185.7,0.0,2570.2,0,0,90277
91,1,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,74.7,74.7,0,79,2,27.65,4182,0,Redondo Beach,0,1,DSL,33.873395,-118.37019,0,74.7,0,0,None,37322,1,0,0,0,1,0,0.0,27.65,0.0,74.7,0,1,90278
92,1,0,1,1,66,1,1,DSL,1,0,1,1,Two year,1,Mailed check,84.0,5714.25,0,57,26,6.22,5825,0,South Gate,1,1,Fiber Optic,33.944624,-118.19261499999999,1,84.0,0,0,Offer A,96267,1,0,0,1,66,1,1486.0,410.52,0.0,5714.25,0,0,90280
93,0,0,0,0,65,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),111.05,7107,0,50,14,41.78,5261,0,Topanga,1,0,DSL,34.115192,-118.61017,0,111.05,0,0,None,5451,0,0,0,1,65,0,995.0,2715.7000000000007,0.0,7107.0,0,0,90290
94,1,0,0,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),100.9,7459.05,0,52,12,24.53,5781,0,Venice,1,1,Fiber Optic,33.991782,-118.479229,0,100.9,0,0,Offer A,31021,0,0,0,1,72,1,895.0,1766.16,0.0,7459.05,0,0,90291
95,0,0,0,0,12,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,78.95,927.35,1,34,62,25.34,5806,1,Marina Del Rey,0,0,DSL,33.977468,-118.445475,0,82.10799999999999,3,0,None,18058,0,0,0,0,12,5,575.0,304.08,0.0,927.35,0,0,90292
96,1,0,1,1,71,1,1,DSL,1,1,0,0,One year,1,Credit card (automatic),66.85,4748.7,0,50,26,4.85,4117,0,Playa Del Rey,0,1,Fiber Optic,33.947305,-118.43984099999999,1,66.85,0,1,Offer A,11264,1,0,1,0,71,0,0.0,344.35,0.0,4748.7,0,1,90293
97,1,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,21.05,113.85,1,30,0,34.26,2604,1,Inglewood,0,1,NA,33.956445,-118.35863400000001,0,21.05,0,0,Offer E,37527,0,1,0,0,5,5,0.0,171.29999999999995,0.0,113.85,0,0,90301
98,1,0,0,0,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),21.0,1107.2,0,62,0,28.3,4158,0,Inglewood,0,1,NA,33.975332,-118.35525200000001,0,21.0,0,0,None,30779,0,0,0,0,52,1,0.0,1471.6,0.0,1107.2,0,0,90302
99,0,1,1,0,25,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,98.5,2514.5,1,78,13,19.76,5337,1,Inglewood,1,0,Fiber Optic,33.936291,-118.33263899999999,1,102.44,1,1,Offer C,27778,0,1,1,0,25,1,327.0,494.00000000000006,13.43,2514.5,0,0,90303
100,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.2,20.2,0,19,0,41.1,2710,0,Inglewood,0,1,NA,33.936827,-118.359824,0,20.2,0,0,Offer E,28680,0,0,0,0,1,3,0.0,41.1,0.0,20.2,1,0,90304
101,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.45,19.45,0,38,0,16.44,5612,0,Inglewood,0,0,NA,33.958134,-118.330905,1,19.45,2,1,Offer E,13779,0,0,1,0,1,1,0.0,16.44,0.0,19.45,0,0,90305
102,1,0,0,0,38,1,1,Fiber optic,0,0,1,0,One year,0,Bank transfer (automatic),95.0,3605.6,0,34,21,3.95,4741,0,Santa Monica,1,1,Fiber Optic,34.015481,-118.49323100000001,0,95.0,0,0,Offer C,5221,1,1,0,0,38,2,75.72,150.1,0.0,3605.6,0,1,90401
103,0,1,1,0,66,0,No phone service,DSL,0,1,1,0,One year,0,Bank transfer (automatic),45.55,3027.25,0,65,9,0.0,6238,0,Santa Monica,1,0,Cable,34.035849,-118.50350800000001,1,45.55,0,0,Offer A,11509,0,0,0,0,66,0,272.0,0.0,0.0,3027.25,0,0,90402
104,1,0,1,0,68,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),110.0,7611.85,1,26,52,14.79,5034,1,Santa Monica,1,1,Cable,34.031529,-118.491156,1,114.4,0,4,Offer A,23559,1,3,1,1,68,1,3958.0,1005.72,0.0,7611.85,1,0,90403
105,1,0,0,0,5,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,24.3,100.2,0,35,21,0.0,4015,0,Santa Monica,0,1,Fiber Optic,34.026334000000006,-118.474222,0,24.3,0,0,Offer E,19975,0,1,0,0,5,1,0.0,0.0,0.0,100.2,0,1,90404
106,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,104.15,7303.05,0,25,59,25.82,4594,0,Santa Monica,0,0,DSL,34.005439,-118.477507,1,104.15,0,1,Offer A,26099,0,0,1,1,72,0,0.0,1859.04,0.0,7303.05,1,1,90405
107,0,0,0,0,32,0,No phone service,DSL,1,0,0,0,One year,0,Mailed check,30.15,927.65,0,60,18,0.0,3585,0,Torrance,0,0,Fiber Optic,33.833698999999996,-118.31438700000001,0,30.15,0,0,Offer C,40705,0,0,0,0,32,1,0.0,0.0,0.0,927.65,0,1,90501
108,1,0,0,0,43,1,1,Fiber optic,0,0,1,1,One year,0,Mailed check,94.35,3921.3,0,50,7,41.22,5845,0,Torrance,0,1,Fiber Optic,33.833181,-118.29206200000002,0,94.35,0,0,None,17058,0,1,0,1,43,3,274.0,1772.46,0.0,3921.3,0,0,90502
109,1,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.4,1363.25,0,38,0,49.5,5234,0,Torrance,0,1,NA,33.840399,-118.353714,1,19.4,0,1,Offer A,41979,0,0,1,0,72,0,0.0,3564.0,0.0,1363.25,0,0,90503
110,1,0,1,0,55,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,96.75,5238.9,1,37,30,49.06,5154,1,Torrance,0,1,DSL,33.867257,-118.330794,1,100.62,1,0,None,31678,0,0,0,0,55,0,1572.0,2698.3,0.0,5238.9,0,0,90504
111,0,0,0,0,52,1,0,DSL,1,0,0,0,One year,0,Credit card (automatic),57.95,3042.25,0,35,5,33.84,6078,0,Torrance,1,0,Cable,33.807882,-118.34795700000001,0,57.95,0,0,None,34873,1,0,0,0,52,1,152.0,1759.6800000000005,0.0,3042.25,0,0,90505
112,0,0,0,0,43,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,91.65,3954.1,0,36,12,26.55,3826,0,Whittier,1,0,Fiber Optic,34.007353,-118.03368300000001,0,91.65,0,0,None,32050,0,0,0,0,43,0,474.0,1141.65,0.0,3954.1,0,0,90601
113,0,1,1,0,37,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.5,2868.15,1,80,15,6.33,2793,1,Whittier,0,0,Cable,33.972119,-118.02018799999999,1,79.56,1,1,Offer C,26265,0,0,1,0,37,1,430.0,234.21,0.0,2868.15,0,0,90602
114,0,0,1,1,64,0,No phone service,DSL,0,1,1,1,Two year,1,Electronic check,54.6,3423.5,0,48,30,0.0,4850,0,Whittier,0,0,DSL,33.945318,-117.992066,1,54.6,0,1,None,19109,1,0,1,1,64,0,1027.0,0.0,0.0,3423.5,0,0,90603
115,1,0,1,1,3,1,0,Fiber optic,1,1,1,0,Month-to-month,0,Electronic check,89.85,248.4,0,38,12,33.3,4648,0,Whittier,0,1,Fiber Optic,33.929704,-118.01208000000001,1,89.85,2,1,Offer E,37887,0,2,1,0,3,1,0.0,99.9,0.0,248.4,0,1,90604
116,0,0,0,0,36,0,No phone service,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),31.05,1126.35,0,61,27,0.0,4871,0,Whittier,0,0,Fiber Optic,33.960891,-118.03222199999999,0,31.05,0,0,Offer C,38181,0,0,0,0,36,3,0.0,0.0,0.0,1126.35,0,1,90605
117,0,0,1,1,10,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,100.25,1064.65,1,62,33,24.48,5998,1,Whittier,0,0,Cable,33.976678,-118.065875,1,104.26,2,1,None,32148,0,2,1,1,10,2,0.0,244.8,0.0,1064.65,0,1,90606
118,0,0,0,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.65,835.15,0,53,0,31.62,5918,0,Buena Park,0,0,NA,33.845706,-118.012204,0,20.65,0,0,None,44442,0,0,0,0,41,1,0.0,1296.42,0.0,835.15,0,0,90620
119,1,0,1,1,27,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),85.2,2151.6,0,33,15,48.17,3796,0,Buena Park,0,1,Fiber Optic,33.874224,-117.99336799999999,1,85.2,1,1,Offer C,33528,1,2,1,0,27,1,323.0,1300.59,0.0,2151.6,0,0,90621
120,0,0,1,1,56,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),99.8,5515.45,0,27,71,42.37,4606,0,La Palma,1,0,DSL,33.850504,-118.039892,1,99.8,0,1,None,15505,0,0,1,1,56,0,0.0,2372.72,0.0,5515.45,1,1,90623
121,0,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.7,112.75,0,31,0,7.72,5346,0,Cypress,0,0,NA,33.818477,-118.038307,0,20.7,0,0,Offer E,47344,0,1,0,0,6,1,0.0,46.32,0.0,112.75,0,0,90630
122,1,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.4,229.55,1,21,78,14.6,4415,1,La Habra,0,1,Cable,33.940619,-117.9513,0,77.376,2,0,Offer E,67354,0,2,0,1,3,3,179.0,43.8,8.74,229.55,1,0,90631
123,0,0,1,1,7,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,50.7,350.35,0,20,71,25.64,3097,0,La Mirada,0,0,Fiber Optic,33.902045,-118.00896100000001,1,50.7,2,1,None,47568,0,2,1,0,7,1,249.0,179.48000000000005,0.0,350.35,1,0,90638
124,0,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.85,62.9,0,27,0,39.89,3172,0,Montebello,0,0,NA,34.015217,-118.10996200000001,1,20.85,1,1,None,62425,0,0,1,0,4,1,0.0,159.56,0.0,62.9,1,0,90640
125,1,0,0,0,33,1,0,Fiber optic,1,0,1,0,Two year,1,Electronic check,88.95,3027.65,0,59,18,47.64,5087,0,Norwalk,0,1,Fiber Optic,33.905963,-118.08263000000001,0,88.95,0,0,Offer C,103214,1,0,0,0,33,0,545.0,1572.12,0.0,3027.65,0,0,90650
126,0,1,0,0,27,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,78.05,2135.5,1,72,20,3.33,4638,1,Pico Rivera,1,0,Fiber Optic,33.989523999999996,-118.089299,0,81.172,1,0,Offer C,63288,0,0,0,0,27,0,427.0,89.91,0.0,2135.5,0,0,90660
127,1,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),23.55,1723.95,0,46,0,1.86,5901,0,Santa Fe Springs,0,1,NA,33.933565,-118.062611,1,23.55,0,1,Offer A,16271,0,0,1,0,72,1,0.0,133.92000000000002,0.0,1723.95,0,0,90670
128,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.75,19.75,0,45,0,15.77,2484,0,Stanton,0,1,NA,33.801869,-117.99506799999999,0,19.75,0,0,None,29694,0,0,0,0,1,2,0.0,15.77,0.0,19.75,0,0,90680
129,1,1,0,0,71,0,No phone service,DSL,1,1,1,1,One year,1,Electronic check,56.45,3985.35,0,73,20,0.0,5372,0,Artesia,0,1,Fiber Optic,33.867593,-118.08063700000001,0,56.45,0,0,Offer A,16398,0,0,0,1,71,2,79.71,0.0,0.0,3985.35,0,1,90701
130,0,0,0,0,13,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.95,1215.65,0,49,22,29.21,5886,0,Cerritos,0,0,DSL,33.8681,-118.067402,0,85.95,0,0,None,51556,0,0,0,1,13,0,26.74,379.73,0.0,1215.65,0,1,90703
131,0,0,1,1,25,0,No phone service,DSL,1,1,1,1,Month-to-month,1,Credit card (automatic),58.6,1502.65,1,27,53,0.0,4190,1,Avalon,1,0,Cable,33.391181,-118.421305,1,60.943999999999996,0,6,Offer C,3699,0,0,1,1,25,3,79.64,0.0,4.48,1502.65,1,1,90704
132,1,0,0,0,67,1,0,DSL,0,0,0,0,Two year,0,Bank transfer (automatic),50.55,3260.1,0,60,8,32.58,6064,0,Bellflower,0,1,DSL,33.887676,-118.12728899999999,0,50.55,0,0,Offer A,72893,1,0,0,0,67,1,0.0,2182.86,0.0,3260.1,0,1,90706
133,1,0,0,0,1,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,35.45,35.45,1,64,24,0.0,2301,1,Harbor City,0,1,Fiber Optic,33.798266,-118.30023700000001,0,36.868,0,0,Offer E,24660,0,1,0,1,1,2,0.0,0.0,0.0,35.45,0,1,90710
134,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.35,81.25,1,45,3,46.84,2570,1,Lakewood,0,1,DSL,33.840524,-118.148403,0,46.123999999999995,0,0,Offer E,30173,0,2,0,0,2,5,2.0,93.68,0.0,81.25,0,0,90712
135,0,0,0,0,43,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.7,1188.2,0,42,0,25.53,2017,0,Lakewood,0,0,NA,33.847755,-118.112532,0,25.7,0,0,None,27563,0,0,0,0,43,0,0.0,1097.79,0.0,1188.2,0,0,90713
136,0,0,0,0,23,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),75.0,1778.5,0,37,22,24.04,2221,0,Lakewood,0,0,Cable,33.841027000000004,-118.078097,0,75.0,0,0,None,20890,0,0,0,0,23,0,391.0,552.92,0.0,1778.5,0,0,90715
137,0,0,1,1,64,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.2,1277.75,0,23,0,36.24,4557,0,Hawaiian Gardens,0,0,NA,33.830431,-118.07407099999999,1,20.2,0,1,None,14852,0,0,1,0,64,0,0.0,2319.36,0.0,1277.75,1,0,90716
138,1,0,0,1,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.6,1170.55,0,58,0,5.71,4393,0,Lomita,0,1,NA,33.794209,-118.31735400000001,0,19.6,0,0,None,21065,0,0,0,0,57,2,0.0,325.47,0.0,1170.55,0,0,90717
139,0,1,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.45,70.45,1,76,33,15.28,3964,1,Los Alamitos,0,0,Cable,33.794990000000006,-118.065591,1,73.268,2,1,Offer E,21343,0,0,1,0,1,7,0.0,15.28,0.0,70.45,0,0,90720
140,0,1,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),88.05,6425.65,0,71,6,20.48,6102,0,Paramount,1,0,Fiber Optic,33.897121999999996,-118.164432,1,88.05,0,1,Offer A,55306,1,0,1,1,72,2,38.55,1474.56,0.0,6425.65,0,1,90723
141,0,0,0,0,8,1,1,DSL,1,0,0,1,Month-to-month,0,Electronic check,71.15,563.65,1,53,20,48.14,2662,1,San Pedro,0,0,DSL,33.736387,-118.28436299999998,0,73.99600000000002,0,0,Offer E,58639,1,0,0,1,8,3,113.0,385.12,0.0,563.65,0,0,90731
142,0,0,1,0,61,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),101.05,5971.25,0,35,21,17.49,6311,0,San Pedro,0,0,Cable,33.744119,-118.31448,1,101.05,0,2,None,21279,0,0,1,1,61,0,0.0,1066.89,0.0,5971.25,0,1,90732
143,1,0,0,0,64,1,1,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),84.3,5289.05,0,34,12,30.27,5044,0,Seal Beach,0,1,DSL,33.75462,-118.071128,0,84.3,0,0,None,24180,0,1,0,0,64,4,635.0,1937.28,0.0,5289.05,0,0,90740
144,1,1,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),23.95,1756.2,0,66,0,30.72,4329,0,Sunset Beach,0,1,NA,33.719221000000005,-118.073596,1,23.95,0,7,Offer A,1107,0,0,1,0,71,1,0.0,2181.12,0.0,1756.2,0,0,90742
145,0,0,1,1,65,1,1,Fiber optic,1,1,1,0,Two year,1,Credit card (automatic),99.05,6416.7,0,56,13,13.2,5878,0,Surfside,0,0,DSL,33.728273,-118.08530400000001,1,99.05,0,5,None,174,1,2,1,0,65,2,83.42,858.0,0.0,6416.7,0,1,90743
146,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.6,61.35,0,42,0,35.65,2543,0,Wilmington,0,1,NA,33.782068,-118.26226299999999,0,19.6,0,0,None,53323,0,0,0,0,3,1,0.0,106.95,0.0,61.35,0,0,90744
147,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.65,45.65,1,63,26,14.12,2600,1,Carson,0,1,DSL,33.822295000000004,-118.26411,0,47.476000000000006,0,0,Offer E,55486,0,2,0,0,1,3,0.0,14.12,0.0,45.65,0,0,90745
148,1,0,0,1,30,1,0,DSL,0,1,1,0,One year,0,Credit card (automatic),64.5,1929.95,0,52,6,27.88,4320,0,Carson,1,1,DSL,33.859171,-118.25227199999999,0,64.5,0,0,Offer C,25566,0,0,0,0,30,1,116.0,836.4,0.0,1929.95,0,0,90746
149,1,0,1,1,15,1,0,DSL,0,1,0,1,Month-to-month,1,Mailed check,69.5,1071.4,0,50,21,8.44,3128,0,Long Beach,1,1,DSL,33.752524,-118.21073700000001,1,69.5,1,1,None,38427,1,1,1,1,15,1,225.0,126.6,0.0,1071.4,0,0,90802
150,0,0,1,1,8,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,68.55,564.35,0,33,17,29.94,3123,0,Long Beach,0,0,Cable,33.760458,-118.129725,1,68.55,1,1,None,31352,1,0,1,1,8,0,96.0,239.52,0.0,564.35,0,0,90803
151,1,0,0,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Mailed check,95.0,655.5,1,32,31,20.52,2786,1,Long Beach,0,1,Cable,33.783046999999996,-118.1486,0,98.8,4,0,Offer E,43467,0,0,0,1,7,0,203.0,143.64,36.6,655.5,0,0,90804
152,0,0,1,1,70,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),108.15,7930.55,0,27,48,5.77,5192,0,Long Beach,1,0,Fiber Optic,33.864622,-118.179626,1,108.15,0,4,Offer A,91664,0,1,1,1,70,1,3807.0,403.9,0.0,7930.55,1,0,90805
153,1,0,1,1,62,1,0,DSL,1,1,1,1,Two year,0,Electronic check,86.1,5215.25,0,51,23,43.2,5769,0,Long Beach,1,1,Cable,33.802664,-118.179971,1,86.1,0,2,None,49647,1,2,1,1,62,1,119.95,2678.4,0.0,5215.25,0,1,90806
154,0,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.7,113.5,0,29,0,5.52,4293,0,Long Beach,0,0,NA,33.830099,-118.182239,1,19.7,3,9,None,31556,0,0,1,0,6,1,0.0,33.12,0.0,113.5,1,0,90807
155,0,0,1,1,14,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),80.9,1152.8,0,33,19,40.22,2563,0,Long Beach,0,0,DSL,33.823943,-118.11133500000001,1,80.9,1,7,None,37417,0,1,1,1,14,1,219.0,563.0799999999998,0.0,1152.8,0,0,90808
156,0,0,0,0,22,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),84.15,1821.95,0,23,41,19.2,3549,0,Long Beach,0,0,Fiber Optic,33.819814,-118.222416,0,84.15,0,0,None,35656,0,0,0,0,22,0,0.0,422.4,0.0,1821.95,1,1,90810
157,1,0,1,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.15,419.9,0,37,0,48.06,2173,0,Long Beach,0,1,NA,33.781086,-118.199049,1,20.15,0,3,None,63136,0,0,1,0,22,2,0.0,1057.3200000000004,0.0,419.9,0,0,90813
158,1,0,1,1,16,1,0,DSL,1,0,1,0,Two year,0,Mailed check,64.25,1024,0,38,27,23.31,5511,0,Long Beach,1,1,Fiber Optic,33.771612,-118.14386599999999,1,64.25,0,9,None,19034,0,0,1,0,16,0,27.65,372.96,0.0,1024.0,0,1,90814
159,1,0,0,0,10,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.7,251.6,0,44,0,32.1,3611,0,Long Beach,0,1,NA,33.797638,-118.11662,0,25.7,0,0,None,38902,0,1,0,0,10,1,0.0,321.0,0.0,251.6,0,0,90815
160,0,0,0,1,13,1,0,DSL,1,1,0,0,Month-to-month,1,Electronic check,56.0,764.55,0,63,10,27.04,5156,0,Long Beach,0,0,Fiber Optic,33.778436,-118.118648,0,56.0,1,0,None,425,0,0,0,0,13,0,7.65,351.52,0.0,764.55,0,1,90822
161,0,0,1,0,20,1,1,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,82.4,1592.35,1,26,56,36.6,5719,1,Altadena,0,0,Fiber Optic,34.196837,-118.14223600000001,1,85.69600000000001,1,5,None,36243,0,1,1,1,20,1,892.0,732.0,33.43,1592.35,1,0,91001
162,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.7,135.2,0,54,8,15.67,3056,0,Arcadia,0,0,Fiber Optic,34.137319,-118.02983700000001,0,69.7,0,0,None,30028,0,0,0,0,2,2,11.0,31.34,0.0,135.2,0,0,91006
163,1,0,0,0,53,1,1,DSL,0,1,0,1,Two year,1,Bank transfer (automatic),73.9,3958.25,0,35,4,6.54,5644,0,Arcadia,1,1,Cable,34.128284,-118.04773200000001,0,73.9,0,0,None,30933,1,0,0,1,53,0,0.0,346.62,0.0,3958.25,0,1,91007
164,0,0,1,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.6,233.9,0,21,0,1.92,4047,0,Duarte,0,0,NA,34.145695,-117.95982,1,20.6,0,7,None,27414,0,0,1,0,11,3,0.0,21.12,0.0,233.9,1,0,91010
165,1,0,1,0,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.9,1363.45,0,40,0,30.86,5570,0,La Canada Flintridge,0,1,NA,34.234912,-118.153729,1,19.9,0,3,Offer A,20200,0,0,1,0,69,0,0.0,2129.34,0.0,1363.45,0,0,91011
166,0,0,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),70.9,273,1,42,30,33.5,4287,1,Monrovia,0,0,Fiber Optic,34.1528,-118.000482,0,73.736,1,0,Offer E,41067,0,3,0,0,4,2,82.0,134.0,8.74,273.0,0,0,91016
167,1,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),89.05,6254.45,0,39,30,6.05,6212,0,Montrose,1,1,DSL,34.2112,-118.230625,1,89.05,0,7,Offer A,7527,1,0,1,1,72,0,0.0,435.6,0.0,6254.45,0,1,91020
168,1,1,1,0,58,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Electronic check,45.3,2651.2,1,66,26,0.0,5444,1,Sierra Madre,1,1,Cable,34.168686,-118.057505,1,47.111999999999995,0,6,Offer B,10558,0,1,1,0,58,2,689.0,0.0,40.95,2651.2,0,0,91024
169,0,0,1,1,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.4,321.4,0,59,0,45.54,3990,0,South Pasadena,0,0,NA,34.110444,-118.156957,1,20.4,2,3,Offer D,23984,0,0,1,0,16,4,0.0,728.64,0.0,321.4,0,0,91030
170,1,0,1,0,43,1,0,Fiber optic,1,0,0,0,One year,1,Bank transfer (automatic),84.25,3539.25,0,61,21,15.2,4382,0,Sunland,1,1,Fiber Optic,34.282703999999995,-118.312929,1,84.25,0,6,None,18752,1,0,1,0,43,3,74.32,653.6,0.0,3539.25,0,1,91040
171,0,0,1,0,2,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,104.4,242.8,1,26,58,11.51,4690,1,Tujunga,1,0,DSL,34.296574,-118.24483899999998,1,108.576,3,1,Offer E,26753,1,2,1,1,2,5,141.0,23.02,45.44,242.8,1,0,91042
172,1,0,1,0,14,1,0,DSL,0,1,1,1,Two year,0,Mailed check,81.95,1181.75,0,48,25,5.17,2564,0,Pasadena,1,1,Cable,34.146634999999996,-118.139225,1,81.95,0,3,Offer D,16812,1,0,1,1,14,1,0.0,72.38,0.0,1181.75,0,1,91101
173,0,0,1,0,53,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),94.85,5000.2,1,24,80,40.62,4328,1,Pasadena,1,0,DSL,34.167465,-118.165327,1,98.644,0,5,None,27891,0,1,1,1,53,3,4000.0,2152.86,18.55,5000.2,1,0,91103
174,0,0,0,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.55,654.55,0,61,0,35.97,5358,0,Pasadena,0,0,NA,34.165383,-118.123752,0,20.55,0,0,Offer C,38460,0,0,0,0,32,2,0.0,1151.04,0.0,654.55,0,0,91104
175,0,0,1,0,34,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,24.7,780.2,0,49,0,11.52,3421,0,Pasadena,0,0,NA,34.13946,-118.16664899999999,1,24.7,0,5,Offer C,10253,0,0,1,0,34,0,0.0,391.68,0.0,780.2,0,0,91105
176,0,1,0,0,15,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.45,1145.7,1,70,21,44.07,5717,1,Pasadena,0,0,Cable,34.139402000000004,-118.128658,0,77.42800000000003,2,0,Offer D,23742,0,0,0,0,15,3,241.0,661.05,0.0,1145.7,0,0,91106
177,0,1,0,0,7,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Bank transfer (automatic),76.45,503.6,1,77,20,26.95,4419,1,Pasadena,0,0,DSL,34.159007,-118.08735300000001,0,79.50800000000002,2,0,Offer E,32369,0,0,0,0,7,3,101.0,188.65,11.05,503.6,0,0,91107
178,0,0,1,1,15,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),105.35,1559.25,0,19,59,4.19,2721,0,San Marino,1,0,Fiber Optic,34.122671000000004,-118.11291100000001,1,105.35,3,6,Offer D,13158,0,0,1,1,15,0,920.0,62.85000000000001,0.0,1559.25,1,0,91108
179,1,0,1,0,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.55,1252,0,22,0,19.27,5110,0,Glendale,0,1,NA,34.17051,-118.28946299999998,1,20.55,0,3,None,23981,0,0,1,0,61,2,0.0,1175.47,0.0,1252.0,1,0,91201
180,0,0,0,0,1,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),29.95,29.95,1,54,30,0.0,4534,1,Glendale,0,0,Cable,34.167926,-118.26753899999999,0,31.148000000000003,0,0,Offer E,21990,0,4,0,0,1,4,0.0,0.0,0.0,29.95,0,0,91202
181,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.3,45.3,0,25,41,47.36,3575,0,Glendale,0,0,Fiber Optic,34.153338,-118.262974,0,45.3,0,0,None,14493,0,0,0,0,1,0,0.0,47.36,0.0,45.3,1,1,91203
182,1,0,0,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Bank transfer (automatic),84.5,662.65,1,51,21,25.73,2152,1,Glendale,0,1,Cable,34.136306,-118.26036,0,87.88000000000002,2,0,Offer E,17015,0,2,0,1,8,4,139.0,205.84,33.21,662.65,0,0,91204
183,1,0,1,1,33,1,0,DSL,1,0,1,1,One year,0,Credit card (automatic),74.75,2453.3,0,35,30,48.85,5344,0,Glendale,1,1,Fiber Optic,34.13658,-118.24583899999999,1,74.75,0,7,Offer C,41390,0,0,1,1,33,3,736.0,1612.05,0.0,2453.3,0,0,91205
184,0,0,0,0,13,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.25,1111.65,1,48,84,33.54,5142,1,Glendale,1,0,DSL,34.162515,-118.203869,0,82.42,3,0,None,31297,0,4,0,0,13,2,934.0,436.02,48.25,1111.65,0,0,91206
185,0,0,1,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.8,24.8,1,29,32,0.0,4851,1,Glendale,0,0,Cable,34.182378,-118.262922,1,25.791999999999998,0,4,Offer E,9864,0,0,1,1,1,0,0.0,0.0,0.0,24.8,1,0,91207
186,1,0,0,0,20,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,51.8,1023.85,0,45,18,3.94,2764,0,Glendale,0,1,DSL,34.195386,-118.23850800000001,0,51.8,0,0,Offer D,16910,0,0,0,0,20,0,184.0,78.8,0.0,1023.85,0,0,91208
187,1,0,0,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,30.4,82.15,0,19,59,0.0,3108,0,La Crescenta,0,1,Cable,34.239636,-118.245259,0,30.4,0,0,None,29110,1,0,0,0,3,1,4.85,0.0,0.0,82.15,1,1,91214
188,0,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.65,244.8,0,61,0,33.13,2024,0,Agoura Hills,0,0,NA,34.129058,-118.75978799999999,0,19.65,0,0,Offer D,25303,0,0,0,0,13,1,0.0,430.69000000000005,0.0,244.8,0,0,91301
189,0,0,1,0,40,1,1,DSL,0,1,0,0,Month-to-month,0,Credit card (automatic),56.6,2379.1,0,62,23,48.29,3359,0,Calabasas,0,0,Fiber Optic,34.130860999999996,-118.68346000000001,1,56.6,0,5,None,23661,0,1,1,0,40,1,0.0,1931.6,0.0,2379.1,0,1,91302
190,1,0,1,1,43,1,1,DSL,1,0,0,1,One year,1,Credit card (automatic),71.9,3173.35,0,24,51,48.1,4106,0,Canoga Park,0,1,Fiber Optic,34.19829,-118.602203,1,71.9,0,5,Offer B,23519,1,0,1,1,43,1,161.84,2068.3,0.0,3173.35,1,1,91303
191,1,0,1,0,6,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,91.0,531,1,39,32,42.08,2283,1,Canoga Park,1,1,Fiber Optic,34.224377000000004,-118.63265600000001,1,94.64,2,5,None,49242,0,1,1,1,6,4,0.0,252.48,0.0,531.0,0,1,91304
192,0,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.75,1375.4,0,38,0,5.27,5325,0,Winnetka,0,0,NA,34.209532,-118.57756299999998,1,19.75,0,9,Offer A,43857,0,0,1,0,69,0,0.0,363.63,0.0,1375.4,0,0,91306
193,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),109.7,8129.3,0,42,3,18.66,5945,0,West Hills,1,0,DSL,34.199787,-118.68493000000001,1,109.7,0,7,Offer A,23637,0,0,1,1,72,2,0.0,1343.52,0.0,8129.3,0,1,91307
194,1,0,1,1,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.3,1192.7,0,33,0,25.57,4149,0,Chatsworth,0,1,NA,34.294142,-118.60388300000001,1,19.3,0,3,Offer B,35325,0,0,1,0,59,2,0.0,1508.63,0.0,1192.7,0,0,91311
195,0,0,1,0,20,1,0,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,96.55,1901.65,0,32,15,28.57,4382,0,Encino,0,0,DSL,34.150354,-118.51829199999999,1,96.55,0,0,Offer D,27614,1,0,0,0,20,0,285.0,571.4,0.0,1901.65,0,0,91316
196,1,0,1,1,24,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.1,587.4,0,19,0,1.14,4634,0,Newbury Park,0,1,NA,34.172071,-118.946262,1,24.1,3,1,Offer C,37779,0,0,1,0,24,1,0.0,27.36,0.0,587.4,1,0,91320
197,1,0,0,0,59,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,111.35,6519.75,0,19,51,48.12,6047,0,Newhall,1,1,Fiber Optic,34.370378,-118.50411799999999,0,111.35,0,0,Offer B,30742,1,0,0,1,59,1,3325.0,2839.08,0.0,6519.75,1,0,91321
198,1,0,1,1,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),112.25,8041.65,0,42,28,11.66,4099,0,Northridge,1,1,DSL,34.238208,-118.55028999999999,1,112.25,3,2,Offer A,25751,1,0,1,1,72,1,0.0,839.52,0.0,8041.65,0,1,91324
199,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.75,20.75,0,29,0,7.57,3358,0,Northridge,0,1,NA,34.236683,-118.51758799999999,0,20.75,1,0,None,32307,0,0,0,0,1,3,0.0,7.57,0.0,20.75,1,0,91325
200,0,0,1,0,27,1,0,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),101.9,2681.15,0,55,27,20.02,3795,0,Porter Ranch,0,0,Fiber Optic,34.281911,-118.55621799999999,1,101.9,0,0,Offer C,28067,1,1,0,1,27,1,0.0,540.54,0.0,2681.15,0,1,91326
201,0,0,0,0,14,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),80.05,1112.3,0,51,21,1.69,4400,0,Pacoima,0,0,Fiber Optic,34.255441999999995,-118.421314,0,80.05,0,0,Offer D,97318,1,0,0,0,14,0,23.36,23.66,0.0,1112.3,0,1,91331
202,1,0,1,1,71,1,1,Fiber optic,1,0,1,1,Two year,0,Electronic check,105.55,7405.5,0,55,53,25.02,5010,0,Reseda,1,1,DSL,34.200175,-118.540958,1,105.55,3,3,Offer A,68018,0,0,1,1,71,2,0.0,1776.42,0.0,7405.5,0,1,91335
203,1,0,0,1,13,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),78.3,1033.95,0,55,22,31.93,5566,0,San Fernando,0,1,DSL,34.286131,-118.435969,0,78.3,3,0,Offer D,33389,0,1,0,0,13,2,22.75,415.09,0.0,1033.95,0,1,91340
204,1,0,0,0,44,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),68.85,2958.95,0,41,28,1.7,2053,0,Sylmar,0,1,Fiber Optic,34.321621,-118.399841,0,68.85,0,0,Offer B,81986,0,0,0,0,44,2,829.0,74.8,0.0,2958.95,0,0,91342
205,0,0,0,0,33,1,0,Fiber optic,0,1,0,0,One year,1,Bank transfer (automatic),79.95,2684.85,0,64,13,42.29,3118,0,North Hills,0,0,Cable,34.238802,-118.48229599999999,0,79.95,0,0,Offer C,57017,1,0,0,0,33,2,0.0,1395.57,0.0,2684.85,0,1,91343
206,1,0,1,1,72,0,No phone service,DSL,1,1,0,1,Two year,1,Credit card (automatic),55.45,4179.2,0,30,47,0.0,4556,0,Granada Hills,1,1,Fiber Optic,34.291273,-118.505104,1,55.45,0,5,Offer A,48867,1,0,1,1,72,0,1964.0,0.0,0.0,4179.2,0,0,91344
207,1,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,79.9,79.9,1,62,23,23.2,3394,1,Mission Hills,0,1,DSL,34.266389000000004,-118.459744,0,83.096,3,0,None,17112,0,0,0,1,1,2,0.0,23.2,0.0,79.9,0,0,91345
208,0,0,0,0,19,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,106.6,1934.45,1,43,21,28.35,3764,1,Santa Clarita,1,0,Fiber Optic,34.502432,-118.41458999999999,0,110.86399999999999,1,0,None,40077,1,2,0,1,19,3,0.0,538.65,21.72,1934.45,0,1,91350
209,1,0,1,0,64,1,0,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),102.45,6654.1,0,22,69,40.49,6398,0,Canyon Country,1,1,Cable,34.422519,-118.420717,1,102.45,0,10,Offer B,59259,1,0,1,1,64,0,4591.0,2591.36,0.0,6654.1,1,0,91351
210,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),46.0,84.5,1,19,45,49.81,2667,1,Sun Valley,0,1,DSL,34.231053,-118.338307,0,47.84,0,0,None,46639,0,0,0,1,2,3,38.0,99.62,0.0,84.5,1,0,91352
211,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,25.25,25.25,0,40,2,0.0,5858,0,Valencia,0,0,Fiber Optic,34.457005,-118.57372600000001,0,25.25,0,0,None,17846,0,0,0,0,1,0,0.0,0.0,0.0,25.25,0,1,91354
212,1,0,0,1,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,1124.2,0,32,0,15.02,5411,0,Valencia,0,1,NA,34.43987,-118.644609,0,19.75,2,0,Offer B,24977,0,0,0,0,61,0,0.0,916.22,0.0,1124.2,0,0,91355
213,0,0,1,1,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,20.0,540.05,0,23,0,27.72,3800,0,Tarzana,0,0,NA,34.157137,-118.548511,1,20.0,0,6,Offer C,27424,0,2,1,0,29,1,0.0,803.88,0.0,540.05,1,0,91356
214,1,1,1,0,23,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,86.8,1975.85,0,66,2,42.59,5788,0,Thousand Oaks,0,1,Fiber Optic,34.214054,-118.88108999999999,1,86.8,0,1,None,42526,0,0,1,1,23,1,40.0,979.57,0.0,1975.85,0,0,91360
215,0,0,1,0,57,0,No phone service,DSL,1,1,1,1,Month-to-month,1,Bank transfer (automatic),58.75,3437.45,0,45,22,0.0,4115,0,Westlake Village,1,0,Fiber Optic,34.130992,-118.894673,1,58.75,0,1,Offer B,18735,0,0,1,1,57,1,0.0,0.0,0.0,3437.45,0,1,91361
216,1,0,1,1,72,0,No phone service,DSL,1,1,0,0,Two year,0,Credit card (automatic),45.25,3139.8,0,46,17,0.0,5041,0,Thousand Oaks,1,1,DSL,34.191842,-118.822796,1,45.25,0,11,Offer A,33057,1,0,1,0,72,1,0.0,0.0,0.0,3139.8,0,1,91362
217,1,0,1,0,66,0,No phone service,DSL,1,1,1,0,Two year,1,Bank transfer (automatic),56.6,3789.2,0,38,29,0.0,5500,0,Woodland Hills,1,1,Fiber Optic,34.153733,-118.59340800000001,1,56.6,0,1,None,25988,1,0,1,0,66,0,1099.0,0.0,0.0,3789.2,0,0,91364
218,1,0,1,1,65,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),84.2,5324.5,0,51,16,41.57,5256,0,Woodland Hills,1,1,Cable,34.178067999999996,-118.61571399999998,1,84.2,0,8,Offer B,36123,1,0,1,1,65,1,852.0,2702.05,0.0,5324.5,0,0,91367
219,0,0,0,0,8,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),80.0,624.6,0,24,73,39.92,2165,0,Oak Park,0,0,Fiber Optic,34.19225,-118.77687399999999,0,80.0,0,0,None,14814,0,0,0,0,8,2,456.0,319.36,0.0,624.6,1,0,91377
220,0,0,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.15,268.35,1,39,19,29.4,2227,1,Stevenson Ranch,0,0,DSL,34.364153,-118.615583,0,72.956,2,0,None,9937,0,0,0,0,4,0,51.0,117.6,21.69,268.35,0,0,91381
221,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.75,1836.9,0,55,0,32.13,4642,0,Castaic,0,0,NA,34.506627,-118.699048,1,24.75,0,3,None,22177,0,0,1,0,71,1,0.0,2281.23,0.0,1836.9,0,0,91384
222,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,20.2,20.2,0,32,0,44.69,4160,0,Van Nuys,0,1,NA,34.178483,-118.43179099999999,1,20.2,0,8,None,40376,0,0,1,0,1,2,0.0,44.69,0.0,20.2,0,0,91401
223,1,0,1,0,4,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.05,179.35,1,50,24,9.67,3394,1,Fallbrook,0,1,Cable,33.362575,-117.299644,1,52.052,0,2,None,42239,1,0,1,0,4,2,43.0,38.68,0.0,179.35,0,0,92028
224,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.35,219.35,0,53,0,16.72,4451,0,Sherman Oaks,0,0,NA,34.147149,-118.463365,0,19.35,0,0,Offer D,22085,0,1,0,0,12,2,0.0,200.64,0.0,219.35,0,0,91403
225,1,0,0,0,24,0,No phone service,DSL,1,0,1,1,One year,1,Mailed check,50.6,1288.75,0,28,46,0.0,4806,0,Van Nuys,0,1,Fiber Optic,34.202494,-118.448048,0,50.6,0,0,Offer C,51348,0,0,0,1,24,1,593.0,0.0,0.0,1288.75,1,0,91405
226,0,0,1,1,31,1,0,DSL,1,0,1,1,One year,1,Mailed check,81.15,2545.75,0,26,41,39.34,5643,0,Van Nuys,1,0,DSL,34.195685,-118.490752,1,81.15,0,2,None,50047,1,1,1,1,31,3,0.0,1219.5400000000004,0.0,2545.75,1,1,91406
227,0,0,1,0,1,1,0,DSL,0,0,1,0,Month-to-month,0,Mailed check,55.2,55.2,1,22,64,35.6,3638,1,Van Nuys,0,0,Fiber Optic,34.178470000000004,-118.45947199999999,1,57.40800000000001,0,0,None,23646,0,0,0,1,1,3,0.0,35.6,0.0,55.2,1,0,91411
228,1,0,0,0,30,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),89.9,2723.15,0,62,2,31.97,3233,0,Sherman Oaks,0,1,Cable,34.146957,-118.432138,0,89.9,0,0,None,29387,1,0,0,1,30,0,54.0,959.1,0.0,2723.15,0,0,91423
229,0,0,1,1,47,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),85.3,4107.25,0,22,52,29.15,5698,0,Encino,0,0,DSL,34.152875,-118.486056,1,85.3,0,6,Offer B,13129,1,0,1,1,47,3,0.0,1370.05,0.0,4107.25,1,1,91436
230,1,0,0,0,54,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),108.0,5760.65,0,49,4,17.76,6370,0,Burbank,0,1,DSL,34.188339,-118.30094199999999,0,108.0,0,0,Offer B,18112,1,0,0,1,54,1,0.0,959.04,0.0,5760.65,0,1,91501
231,1,0,0,0,50,1,0,Fiber optic,1,1,0,1,Month-to-month,1,Credit card (automatic),93.5,4747.5,0,64,21,40.83,6367,0,Burbank,0,1,DSL,34.177267,-118.31003,0,93.5,0,0,Offer B,11517,1,0,0,1,50,0,0.0,2041.5,0.0,4747.5,0,1,91502
232,1,0,0,0,1,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Mailed check,84.6,84.6,1,40,12,26.85,2484,1,Burbank,0,1,Fiber Optic,34.213049,-118.317651,0,87.984,1,0,None,25882,0,2,0,1,1,2,0.0,26.85,0.0,84.6,0,1,91504
233,0,0,0,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.25,1566.9,0,62,0,42.36,5733,0,Burbank,0,0,NA,34.174215000000004,-118.345928,0,20.25,0,0,None,29245,0,0,0,0,72,0,0.0,3049.92,0.0,1566.9,0,0,91505
234,0,0,0,0,29,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,25.15,702,0,47,0,4.53,5491,0,Burbank,0,0,NA,34.169706,-118.323548,0,25.15,0,0,None,18539,0,0,0,0,29,1,0.0,131.37,0.0,702.0,0,0,91506
235,1,0,0,0,2,1,1,DSL,0,1,0,0,Month-to-month,1,Mailed check,54.4,114.1,1,22,80,44.31,2556,1,North Hollywood,0,1,DSL,34.1692,-118.372498,0,56.576,0,0,None,36625,0,0,0,1,2,0,91.0,88.62,0.0,114.1,1,0,91601
236,0,0,0,0,10,0,No phone service,DSL,0,0,0,0,Two year,1,Mailed check,29.6,299.05,0,41,29,0.0,3180,0,North Hollywood,0,0,Fiber Optic,34.15136,-118.36478600000001,0,29.6,0,0,Offer D,16996,1,2,0,0,10,1,87.0,0.0,0.0,299.05,0,0,91602
237,1,0,1,0,18,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.15,1305.95,0,42,23,16.78,4283,0,Studio City,0,1,Cable,34.139082,-118.39275,1,73.15,0,5,Offer D,26157,0,0,1,0,18,3,30.04,302.04,0.0,1305.95,0,1,91604
238,0,1,0,0,11,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,95.0,1120.3,1,78,32,11.59,5980,1,North Hollywood,0,0,DSL,34.207295,-118.40002199999999,0,98.8,1,0,Offer D,57146,0,2,0,0,11,2,358.0,127.49,0.0,1120.3,0,0,91605
239,1,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,284.35,0,40,0,40.17,4272,0,North Hollywood,0,1,NA,34.187599,-118.387125,0,19.75,0,0,Offer D,45358,0,0,0,0,16,0,0.0,642.72,0.0,284.35,0,0,91606
240,0,0,0,0,72,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),86.6,6350.5,0,37,13,8.29,4530,0,Valley Village,1,0,Cable,34.165783000000005,-118.399795,0,86.6,0,0,None,27453,1,0,0,1,72,1,0.0,596.8799999999999,0.0,6350.5,0,1,91607
241,1,0,0,0,72,1,1,Fiber optic,0,1,1,1,Two year,0,Bank transfer (automatic),109.2,7878.3,0,49,22,35.11,4551,0,Rancho Cucamonga,1,1,Fiber Optic,34.132275,-117.611478,0,109.2,0,0,None,39064,1,0,0,1,72,1,0.0,2527.92,0.0,7878.3,0,1,91701
242,0,0,1,1,41,1,0,DSL,1,0,1,1,One year,1,Credit card (automatic),74.7,3187.65,0,38,11,25.16,5246,0,Azusa,0,0,Cable,34.174493,-117.87068000000001,1,74.7,0,10,Offer B,57775,1,0,1,1,41,1,0.0,1031.56,0.0,3187.65,0,1,91702
243,0,1,1,0,65,1,0,Fiber optic,1,1,0,1,Month-to-month,0,Electronic check,94.4,6126.15,0,77,25,38.32,5348,0,Baldwin Park,1,0,Fiber Optic,34.098275,-117.967399,1,94.4,0,2,None,76890,0,0,1,1,65,0,1532.0,2490.8,0.0,6126.15,0,0,91706
244,0,1,0,0,13,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,54.8,731.3,0,68,20,10.51,5557,0,Chino Hills,1,0,Fiber Optic,33.942895,-117.72564399999999,0,54.8,0,0,None,66754,0,1,0,0,13,1,14.63,136.63,0.0,731.3,0,1,91709
245,1,1,0,0,4,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,75.35,273.4,0,66,29,36.4,4033,0,Chino,0,1,Fiber Optic,33.990646000000005,-117.663025,0,75.35,0,0,Offer E,75319,0,0,0,0,4,0,0.0,145.6,0.0,273.4,0,1,91710
246,1,0,0,0,41,1,1,DSL,0,0,0,1,One year,0,Mailed check,65.0,2531.8,0,35,30,37.55,5043,0,Claremont,1,1,DSL,34.127621000000005,-117.717863,0,65.0,0,0,Offer B,34716,0,0,0,1,41,1,0.0,1539.55,0.0,2531.8,0,1,91711
247,1,1,0,0,15,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.4,1074.3,1,65,32,29.11,4616,1,Covina,0,1,DSL,34.097345000000004,-117.90673600000001,0,77.376,0,0,Offer D,33817,0,0,0,0,15,0,344.0,436.65,0.0,1074.3,0,0,91722
248,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,48.55,48.55,1,37,10,11.35,5687,1,Covina,0,1,Cable,34.084747,-117.886844,0,50.492,0,0,None,17554,0,0,0,0,1,5,0.0,11.35,0.0,48.55,0,0,91723
249,1,0,0,0,42,1,1,Fiber optic,1,1,0,1,One year,1,Electronic check,99.0,4298.45,0,28,48,6.42,2887,0,Covina,1,1,DSL,34.081109999999995,-117.853935,0,99.0,0,0,Offer B,25068,0,0,0,1,42,1,2063.0,269.64,0.0,4298.45,1,0,91724
250,0,0,1,0,51,1,0,Fiber optic,1,1,1,0,One year,1,Electronic check,93.5,4619.55,0,27,46,21.07,5561,0,Rancho Cucamonga,1,0,Fiber Optic,34.100970000000004,-117.57882,1,93.5,0,2,Offer B,51970,0,0,1,0,51,1,0.0,1074.57,0.0,4619.55,1,1,91730
251,0,0,1,1,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.4,147.15,1,47,23,46.23,5687,1,El Monte,0,0,Cable,34.079934,-118.046695,1,73.21600000000002,0,1,None,30211,0,1,1,0,2,1,34.0,92.46,0.0,147.15,0,0,91731
252,1,1,1,0,1,0,No phone service,DSL,0,1,1,0,Month-to-month,0,Electronic check,40.2,40.2,1,77,13,0.0,5828,1,El Monte,0,1,Cable,34.074492,-118.01462,1,41.80800000000001,0,1,Offer E,62660,0,0,1,0,1,2,0.0,0.0,0.0,40.2,0,1,91732
253,1,0,0,1,32,1,1,DSL,0,1,1,1,One year,0,Credit card (automatic),83.7,2633.3,0,56,15,37.48,3945,0,South El Monte,1,1,Fiber Optic,34.04622,-118.053753,0,83.7,0,0,None,45645,1,0,0,1,32,0,0.0,1199.36,0.0,2633.3,0,1,91733
254,1,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.85,193.05,0,29,0,1.98,3768,0,Rancho Cucamonga,0,1,NA,34.245289,-117.642503,0,19.85,0,0,Offer D,23079,0,0,0,0,10,0,0.0,19.8,0.0,193.05,1,0,91737
255,0,0,1,1,67,0,No phone service,DSL,0,1,1,1,Two year,1,Electronic check,59.55,4103.9,0,19,52,0.0,4478,0,Rancho Cucamonga,1,0,Fiber Optic,34.133809,-117.523724,1,59.55,0,1,None,12937,1,0,1,1,67,0,0.0,0.0,0.0,4103.9,1,1,91739
256,0,0,1,1,61,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),115.1,7008.15,0,42,12,20.01,6090,0,Glendora,1,0,Fiber Optic,34.119363,-117.85505900000001,1,115.1,1,3,Offer B,25135,1,0,1,1,61,1,841.0,1220.61,0.0,7008.15,0,0,91740
257,1,0,0,0,50,1,1,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),114.35,5791.1,0,46,21,19.8,5068,0,Glendora,1,1,DSL,34.14649,-117.84981499999999,0,114.35,0,0,Offer B,24973,1,0,0,1,50,2,1216.0,990.0,0.0,5791.1,0,0,91741
258,0,0,1,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),44.6,80.55,1,41,18,30.19,4884,1,La Puente,0,0,DSL,34.031441,-117.93643600000001,1,46.38399999999999,0,3,Offer E,84965,0,0,1,0,2,3,14.0,60.38,0.0,80.55,0,0,91744
259,0,1,1,0,29,0,No phone service,DSL,1,0,0,1,Month-to-month,1,Electronic check,45.0,1228.65,0,69,23,0.0,3094,0,Hacienda Heights,1,0,Fiber Optic,33.998471,-117.973758,1,45.0,0,5,None,53686,0,0,1,0,29,0,0.0,0.0,0.0,1228.65,0,1,91745
260,1,1,0,0,3,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,41.15,132.2,1,67,31,0.0,2314,1,La Puente,1,1,DSL,34.038983,-117.991372,0,42.79600000000001,0,0,Offer E,30802,0,1,0,1,3,7,41.0,0.0,0.0,132.2,0,0,91746
261,1,1,0,0,13,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.9,1364.3,1,68,12,32.68,2494,1,Rowland Heights,1,1,Cable,33.976753,-117.89736699999999,0,111.17600000000002,0,0,Offer D,46342,0,2,0,0,13,1,164.0,424.84,0.0,1364.3,0,0,91748
262,1,1,1,0,57,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.85,4925.35,0,79,9,36.66,4429,0,La Verne,0,1,Cable,34.144703,-117.770299,1,89.85,0,1,None,35530,0,0,1,0,57,0,0.0,2089.62,0.0,4925.35,0,1,91750
263,0,0,0,0,31,0,No phone service,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),49.85,1520.1,0,35,10,0.0,2539,0,Mira Loma,0,0,Fiber Optic,33.999992,-117.535395,0,49.85,0,0,None,18980,1,0,0,1,31,0,0.0,0.0,0.0,1520.1,0,1,91752
264,0,0,1,0,45,1,1,Fiber optic,1,1,1,1,One year,0,Mailed check,113.3,5032.25,0,57,4,33.54,4885,0,Monterey Park,1,0,Fiber Optic,34.050321999999994,-118.14703700000001,1,113.3,0,1,Offer B,33280,1,0,1,1,45,0,0.0,1509.3,0.0,5032.25,0,1,91754
265,0,0,1,1,61,1,1,DSL,1,1,1,1,Two year,0,Mailed check,88.1,5526.75,0,62,28,47.19,5152,0,Monterey Park,1,0,Cable,34.049172,-118.115022,1,88.1,0,1,Offer B,26933,1,0,1,1,61,1,154.75,2878.59,0.0,5526.75,0,1,91755
266,1,0,0,0,50,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.9,1195.25,0,64,0,47.16,4297,0,Mt Baldy,0,1,NA,34.231318,-117.66203200000001,0,24.9,0,0,Offer B,47,0,0,0,0,50,1,0.0,2358.0,0.0,1195.25,0,0,91759
267,0,1,0,0,19,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Mailed check,105.0,2007.25,0,67,12,7.95,3524,0,Ontario,0,0,Fiber Optic,34.035602000000004,-117.591528,0,105.0,0,0,None,56280,1,0,0,0,19,1,24.09,151.05,0.0,2007.25,0,1,91761
268,1,0,0,0,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.35,1099.6,1,51,0,26.63,5084,1,Ontario,0,1,NA,34.057256,-117.667677,0,19.35,0,0,None,54254,0,0,0,0,59,2,0.0,1571.1699999999996,14.22,1099.6,0,0,91762
269,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.25,1732.95,0,30,0,8.21,5409,0,Montclair,0,0,NA,34.072121,-117.698319,1,24.25,0,1,None,34447,0,0,1,0,71,1,0.0,582.9100000000002,0.0,1732.95,0,0,91763
270,0,1,0,0,16,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.45,1511.2,1,68,10,9.43,3810,1,Ontario,0,0,Fiber Optic,34.074087,-117.60561799999999,0,98.228,0,0,Offer D,49474,1,0,0,1,16,0,151.0,150.88,0.0,1511.2,0,0,91764
271,1,0,1,0,57,1,0,DSL,1,1,0,0,Two year,1,Electronic check,59.75,3450.15,0,50,22,49.29,4012,0,Diamond Bar,0,1,Fiber Optic,33.992416,-117.807874,1,59.75,0,1,Offer B,46532,1,0,1,0,57,1,0.0,2809.53,0.0,3450.15,0,1,91765
272,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),24.8,24.8,1,60,32,0.0,5087,1,Pomona,0,1,DSL,34.042286,-117.756106,0,25.791999999999998,0,0,Offer E,69974,0,2,0,0,1,2,0.0,0.0,0.0,24.8,0,0,91766
273,1,1,1,0,20,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,107.05,2172.05,0,68,3,27.56,5328,0,Pomona,0,1,Cable,34.083086,-117.737997,1,107.05,0,3,None,46626,1,0,1,0,20,0,0.0,551.1999999999998,0.0,2172.05,0,1,91767
274,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.6,70.6,1,30,45,44.59,3338,1,Pomona,0,1,Cable,34.067932,-117.785168,0,73.42399999999998,0,0,Offer E,36057,0,0,0,0,1,5,0.0,44.59,0.0,70.6,0,0,91768
275,1,0,1,0,5,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,85.4,401.1,1,51,18,42.29,3676,1,Rosemead,0,1,Fiber Optic,34.065108,-118.08279099999999,1,88.816,0,1,Offer E,61623,1,3,1,0,5,2,72.0,211.45,45.37,401.1,0,0,91770
276,0,0,1,0,52,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.05,5624.85,1,20,53,10.59,4839,1,San Dimas,1,0,DSL,34.102119,-117.815532,1,109.25200000000001,0,6,None,33878,0,0,1,1,52,0,2981.0,550.68,27.6,5624.85,1,0,91773
277,1,1,1,0,21,1,0,DSL,1,1,0,1,Month-to-month,1,Bank transfer (automatic),64.95,1339.8,0,79,30,42.95,4604,0,San Gabriel,0,1,Cable,34.114771999999995,-118.089431,1,64.95,0,5,None,23444,0,0,1,0,21,2,0.0,901.95,0.0,1339.8,0,1,91775
278,1,0,0,0,14,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,55.0,771.95,0,47,4,0.0,4900,0,San Gabriel,1,1,Fiber Optic,34.089927,-118.09564499999999,0,55.0,0,0,Offer D,38041,1,0,0,1,14,2,0.0,0.0,0.0,771.95,0,1,91776
279,0,0,0,0,5,1,0,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),50.55,244.75,0,24,42,43.02,2739,0,Temple City,0,0,Fiber Optic,34.101608,-118.055848,0,50.55,0,0,None,32718,0,0,0,0,5,1,103.0,215.1,0.0,244.75,1,0,91780
280,0,0,0,0,6,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,55.15,322.9,0,29,30,6.98,5377,0,Upland,0,0,Fiber Optic,34.141146,-117.65558300000001,0,55.15,0,0,Offer E,23331,0,0,0,0,6,0,9.69,41.88,0.0,322.9,1,1,91784
281,0,0,0,0,10,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,51.2,498.25,0,44,17,45.56,5765,0,Upland,0,0,Fiber Optic,34.105493,-117.66093400000001,0,51.2,0,0,Offer D,48827,0,1,0,0,10,3,0.0,455.6,0.0,498.25,0,1,91786
282,0,0,0,1,1,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,25.4,25.4,0,21,0,32.73,4556,0,Walnut,0,0,NA,34.018353999999995,-117.85491999999999,0,25.4,1,0,Offer E,45118,0,0,0,0,1,1,0.0,32.73,0.0,25.4,1,0,91789
283,0,0,0,0,68,1,1,DSL,1,0,0,0,Month-to-month,0,Mailed check,54.45,3687.75,0,24,59,5.3,5310,0,West Covina,0,0,Cable,34.066964,-117.93700700000001,0,54.45,0,0,None,44099,0,0,0,0,68,0,2176.0,360.4,0.0,3687.75,1,0,91790
284,1,0,1,1,18,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Mailed check,95.15,1779.95,1,52,31,1.51,4643,1,West Covina,1,1,Fiber Optic,34.061634000000005,-117.893169,1,98.956,0,6,None,30458,0,1,1,1,18,4,552.0,27.18,10.17,1779.95,0,0,91791
285,0,0,0,0,22,1,1,Fiber optic,0,0,0,0,One year,1,Credit card (automatic),76.0,1783.6,0,64,5,19.72,2031,0,West Covina,0,0,DSL,34.024405,-117.89872199999999,0,76.0,0,0,Offer D,31622,0,0,0,0,22,1,0.0,433.84,0.0,1783.6,0,1,91792
286,0,0,0,0,20,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.35,927.15,0,35,18,4.15,3460,0,Alhambra,0,0,DSL,34.090925,-118.12816399999998,0,44.35,0,0,Offer D,54382,0,0,0,0,20,1,167.0,83.0,0.0,927.15,0,0,91801
287,1,0,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.0,70,1,41,20,19.15,4094,1,Alhambra,0,1,Cable,34.074736,-118.145959,1,72.8,0,1,Offer E,30635,0,0,1,0,1,0,0.0,19.15,0.0,70.0,0,1,91803
288,1,1,0,0,8,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.5,606.55,1,66,8,1.78,4345,1,Alpine,0,1,Cable,32.827184,-116.70372900000001,0,77.48,0,0,None,16486,0,2,0,0,8,5,0.0,14.24,0.0,606.55,0,1,91901
289,1,0,0,0,10,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),44.85,435.4,1,34,19,49.58,4061,1,San Diego,0,1,Fiber Optic,32.85723,-117.209774,0,46.64400000000001,0,0,None,34902,0,0,0,0,10,2,83.0,495.8,0.0,435.4,0,0,92122
290,1,1,0,0,24,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.1,1712.7,1,69,16,30.87,2018,1,San Diego,0,1,Fiber Optic,32.85723,-117.209774,0,79.14399999999998,0,0,Offer C,34902,0,0,0,0,24,0,0.0,740.88,0.0,1712.7,0,1,92122
291,1,0,0,0,35,1,0,DSL,1,1,0,0,One year,0,Mailed check,61.2,2021.2,0,24,82,38.38,2075,0,Campo,1,1,Fiber Optic,32.673483000000004,-116.47286299999999,0,61.2,0,0,None,3133,0,0,0,0,35,3,0.0,1343.3000000000004,0.0,2021.2,1,1,91906
292,1,0,1,1,23,1,0,Fiber optic,0,1,0,0,One year,0,Mailed check,86.8,1940.8,0,51,22,16.63,3200,0,Chula Vista,1,1,Fiber Optic,32.636792,-117.05498899999999,1,86.8,0,2,Offer D,74025,1,0,1,0,23,0,0.0,382.49,0.0,1940.8,0,1,91910
293,0,1,0,0,6,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.35,567.8,0,77,19,8.06,2578,0,Chula Vista,0,0,Fiber Optic,32.607964,-117.059459,0,89.35,0,0,Offer E,71126,0,1,0,0,6,2,0.0,48.36,0.0,567.8,0,1,91911
294,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.7,220.35,0,43,0,18.71,5715,0,Chula Vista,0,0,NA,32.64164,-116.985026,0,19.7,0,0,None,12884,0,0,0,0,12,0,0.0,224.52,0.0,220.35,0,0,91913
295,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,20.25,0,44,0,40.46,5384,0,Chula Vista,0,1,NA,32.688506,-116.93863200000001,0,20.25,0,0,Offer E,2606,0,0,0,0,1,0,0.0,40.46,0.0,20.25,0,0,91914
296,0,0,1,1,71,1,0,Fiber optic,0,0,0,0,Two year,0,Electronic check,76.05,5436.45,0,38,10,9.4,5841,0,Chula Vista,1,0,Fiber Optic,32.605012,-116.97595,1,76.05,1,6,None,9278,0,0,1,0,71,0,0.0,667.4,0.0,5436.45,0,1,91915
297,1,1,1,0,35,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.8,3437.5,0,73,3,2.12,3318,0,Descanso,1,1,DSL,32.912664,-116.63538700000001,1,100.8,0,4,None,1587,0,0,1,0,35,0,0.0,74.2,0.0,3437.5,0,1,91916
298,1,0,1,1,40,1,1,DSL,0,0,1,1,Month-to-month,1,Electronic check,74.55,3015.75,0,32,75,13.86,3718,0,Dulzura,1,1,Fiber Optic,32.622999,-116.687855,1,74.55,3,5,Offer B,727,0,0,1,1,40,2,2262.0,554.4,0.0,3015.75,0,0,91917
299,0,0,0,1,1,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,73.6,73.6,1,21,57,6.19,2565,1,San Diego,0,0,Fiber Optic,32.85723,-117.209774,0,76.544,0,0,None,34902,0,1,0,1,1,4,0.0,6.19,0.0,73.6,1,1,92122
300,1,0,0,0,23,1,0,DSL,0,0,1,1,One year,1,Bank transfer (automatic),64.9,1509.8,0,34,23,46.4,3314,0,Imperial Beach,0,1,DSL,32.579134,-117.119009,0,64.9,0,0,None,26662,0,2,0,1,23,2,34.73,1067.2,0.0,1509.8,0,1,91932
301,0,1,0,0,4,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.45,396.1,1,74,2,31.61,3677,1,San Diego,0,0,Cable,32.85723,-117.209774,0,99.26799999999999,0,0,Offer E,34902,0,0,0,0,4,4,8.0,126.44,0.0,396.1,0,0,92122
302,1,0,0,0,4,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,90.4,356.65,0,55,4,31.92,3314,0,Jamul,1,1,Fiber Optic,32.695681,-116.79838600000001,0,90.4,0,0,None,8759,1,0,0,1,4,0,0.0,127.68,0.0,356.65,0,1,91935
303,0,0,1,1,68,0,No phone service,DSL,0,1,1,1,Two year,0,Credit card (automatic),60.3,4109,0,44,15,0.0,4864,0,La Mesa,1,0,Cable,32.759327,-116.99726000000001,1,60.3,0,8,None,44652,1,0,1,1,68,0,61.64,0.0,0.0,4109.0,0,1,91941
304,1,0,0,1,38,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,81.85,3141.7,0,44,13,1.27,3571,0,La Mesa,0,1,Cable,32.782501,-117.01611000000001,0,81.85,2,0,None,24005,0,0,0,0,38,0,0.0,48.26,0.0,3141.7,0,1,91942
305,1,0,1,1,52,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.8,1229.1,0,42,0,40.33,5320,0,Lemon Grove,0,1,NA,32.733564,-117.03371299999999,1,24.8,3,1,Offer B,24961,0,0,1,0,52,1,0.0,2097.16,0.0,1229.1,0,0,91945
306,1,1,1,0,32,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.9,2303.35,1,76,11,47.34,4105,1,San Diego,0,1,DSL,32.85723,-117.209774,1,77.89600000000002,0,2,Offer C,34902,0,0,1,0,32,4,253.0,1514.88,0.0,2303.35,0,0,92122
307,1,0,1,1,29,1,0,DSL,0,0,1,1,Two year,0,Mailed check,75.55,2054.4,0,60,7,32.46,5625,0,National City,1,1,DSL,32.67102,-117.095235,1,75.55,0,7,None,62355,1,1,1,1,29,2,14.38,941.34,0.0,2054.4,0,1,91950
308,1,1,1,1,38,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,101.15,3741.85,0,71,27,28.3,4036,0,Pine Valley,0,1,DSL,32.800671,-116.48336299999998,1,101.15,1,9,None,1604,0,0,1,0,38,2,0.0,1075.4,0.0,3741.85,0,1,91962
309,1,0,0,1,48,1,1,DSL,1,0,1,1,One year,1,Credit card (automatic),78.75,3682.45,0,51,6,2.53,2257,0,Potrero,1,1,DSL,32.619465000000005,-116.59360500000001,0,78.75,0,0,Offer B,905,0,0,0,1,48,3,22.09,121.44,0.0,3682.45,0,1,91963
310,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.25,19.25,0,34,0,9.44,4745,0,Spring Valley,0,0,NA,32.726627,-116.99460800000001,0,19.25,0,0,Offer E,56100,0,0,0,0,1,2,0.0,9.44,0.0,19.25,0,0,91977
311,0,0,0,0,22,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,89.05,1886.25,0,40,8,6.0,5479,0,Spring Valley,0,0,Fiber Optic,32.730264,-116.95096299999999,0,89.05,0,0,None,7863,1,1,0,1,22,1,0.0,132.0,0.0,1886.25,0,1,91978
312,0,0,0,0,43,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),115.05,4895.1,0,25,26,24.85,4115,0,Tecate,1,0,Fiber Optic,32.587557000000004,-116.636816,0,115.05,0,0,Offer B,91,1,0,0,1,43,1,0.0,1068.55,10.76,4895.1,1,1,91980
313,0,1,1,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.35,341.6,0,67,13,9.56,5437,0,Bonsall,0,0,DSL,33.290907000000004,-117.202895,1,69.35,0,0,Offer E,3849,0,1,0,0,5,1,44.0,47.8,0.0,341.6,0,0,92003
314,1,0,0,0,5,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.6,415.55,1,30,57,5.78,5715,1,San Diego,0,1,DSL,32.85723,-117.209774,0,83.824,0,0,Offer E,34902,0,0,0,0,5,2,0.0,28.9,36.44,415.55,0,1,92122
315,1,0,1,1,51,1,1,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),110.05,5686.4,0,23,41,26.73,5604,0,Cardiff By The Sea,0,1,Fiber Optic,33.015865999999995,-117.272254,1,110.05,0,6,None,10375,1,0,1,1,51,0,233.14,1363.23,20.28,5686.4,1,1,92007
316,1,0,0,0,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.9,1355.1,0,49,0,22.22,5308,0,Carlsbad,0,1,NA,33.148115999999995,-117.30604299999999,0,19.9,0,0,None,35582,0,0,0,0,71,0,0.0,1577.62,42.18,1355.1,0,0,92008
317,0,0,1,1,38,1,0,DSL,1,1,1,1,One year,0,Credit card (automatic),80.3,3058.65,1,55,21,42.14,2071,1,San Diego,0,0,DSL,32.85723,-117.209774,1,83.512,0,1,Offer C,34902,1,1,1,1,38,5,642.0,1601.32,0.0,3058.65,0,0,92122
318,1,1,1,0,24,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.15,2231.05,1,77,13,16.1,2212,1,San Diego,1,1,Fiber Optic,32.85723,-117.209774,1,96.876,0,1,Offer C,34902,0,0,1,1,24,1,0.0,386.4,0.0,2231.05,0,1,92122
319,1,0,1,0,35,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),91.5,3236.35,0,64,10,23.85,3617,0,El Cajon,0,1,Fiber Optic,32.785165,-116.862648,1,91.5,0,2,None,40995,1,0,1,0,35,3,0.0,834.75,40.79,3236.35,0,1,92019
320,0,1,0,0,54,1,1,DSL,1,1,1,1,One year,0,Bank transfer (automatic),82.45,4350.1,1,70,6,12.08,4149,1,San Diego,0,0,DSL,32.85723,-117.209774,0,85.74799999999999,0,0,Offer B,34902,1,0,0,1,54,3,0.0,652.32,0.0,4350.1,0,1,92122
321,0,0,1,1,72,0,No phone service,DSL,0,1,1,1,Two year,1,Electronic check,60.0,4264,0,63,16,0.0,5471,0,El Cajon,1,0,Cable,32.832706,-116.873258,1,60.0,0,3,None,61872,1,0,1,1,72,0,68.22,0.0,25.67,4264.0,0,1,92021
322,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.8,44.8,0,40,26,27.46,2269,0,Encinitas,0,1,DSL,33.054579,-117.25665,0,44.8,0,0,Offer E,47126,0,2,0,0,1,2,0.0,27.46,0.0,44.8,0,1,92024
323,0,0,1,1,9,1,0,DSL,1,0,0,0,One year,0,Mailed check,48.6,422.3,0,31,30,30.07,4562,0,Escondido,0,0,Cable,33.081478000000004,-117.03381399999999,1,48.6,0,9,Offer E,49281,0,0,1,0,9,0,127.0,270.63,20.45,422.3,0,0,92025
324,1,0,0,0,69,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),60.05,4176.7,0,62,18,0.0,5388,0,Escondido,0,1,Fiber Optic,33.21846,-117.11691599999999,0,60.05,0,0,None,43436,1,0,0,1,69,0,75.18,0.0,41.21,4176.7,0,1,92026
325,0,0,1,0,52,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),102.7,5138.1,0,30,71,44.34,4044,0,Escondido,0,0,DSL,33.141265000000004,-116.967221,1,102.7,0,0,None,48690,1,0,0,1,52,2,0.0,2305.6800000000007,0.0,5138.1,0,1,92027
326,0,1,1,0,11,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,82.9,880.05,0,68,2,29.15,4413,0,Fallbrook,0,0,Fiber Optic,33.362575,-117.299644,1,82.9,0,9,Offer D,42239,1,0,1,0,11,3,0.0,320.65,0.0,880.05,0,1,92028
327,0,1,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.35,139.05,1,74,11,13.17,2671,1,San Diego,0,0,Fiber Optic,32.85723,-117.209774,0,73.164,0,0,Offer E,34902,0,0,0,0,2,4,15.0,26.34,0.0,139.05,0,0,92122
328,0,1,1,1,28,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,35.9,973.65,0,75,58,0.0,5444,0,Julian,0,0,Fiber Optic,32.980678000000005,-116.262854,1,35.9,3,3,None,3577,0,0,1,0,28,0,565.0,0.0,0.0,973.65,0,0,92036
329,0,1,0,0,17,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),82.65,1470.05,0,79,25,1.06,3754,0,La Jolla,1,0,Fiber Optic,32.853743,-117.25034,0,82.65,0,0,Offer D,42617,0,0,0,0,17,2,368.0,18.02,0.0,1470.05,0,0,92037
330,0,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.85,739.35,0,37,0,9.04,4177,0,Lakeside,0,0,NA,32.909873,-116.906774,1,19.85,1,5,None,42277,0,0,1,0,35,1,0.0,316.4,2.29,739.35,0,0,92040
331,0,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.2,161.95,0,31,0,31.02,5272,0,Oceanside,0,0,NA,33.351059,-117.420557,0,19.2,0,0,Offer E,98239,0,0,0,0,8,0,0.0,248.16,0.0,161.95,0,0,92054
332,1,0,0,0,46,1,1,Fiber optic,0,1,1,0,One year,1,Credit card (automatic),94.9,4422.95,0,31,22,22.13,5316,0,Oceanside,1,1,Fiber Optic,33.194742,-117.29032,0,94.9,0,0,None,52895,0,0,0,0,46,0,973.0,1017.98,24.08,4422.95,0,0,92056
333,0,0,0,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.85,511.25,1,29,29,28.62,2473,1,San Diego,0,0,Cable,32.85723,-117.209774,0,76.804,0,0,None,34902,0,0,0,1,7,1,148.0,200.34,13.03,511.25,1,0,92122
334,0,0,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,80.6,155.8,1,54,22,5.32,2683,1,San Diego,1,0,Cable,32.85723,-117.209774,0,83.824,0,0,None,34902,0,1,0,0,2,3,34.0,10.64,0.0,155.8,0,0,92122
335,1,0,1,1,68,1,1,DSL,0,1,0,1,One year,1,Bank transfer (automatic),75.8,5293.95,1,63,20,29.18,4903,1,San Diego,1,1,Fiber Optic,32.85723,-117.209774,1,78.832,0,1,Offer A,34902,1,0,1,1,68,0,1059.0,1984.24,0.0,5293.95,0,0,92122
336,0,0,0,0,43,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,104.6,4759.85,1,24,65,12.88,5250,1,San Diego,1,0,Fiber Optic,32.85723,-117.209774,0,108.784,0,0,None,34902,0,0,0,1,43,1,0.0,553.84,0.0,4759.85,1,1,92122
337,0,0,0,0,68,1,1,DSL,1,1,1,1,Two year,1,Electronic check,88.15,6148.45,0,63,2,21.82,5531,0,Poway,1,0,Fiber Optic,32.984395,-117.01345400000001,0,88.15,0,0,None,47969,1,0,0,1,68,0,123.0,1483.76,36.29,6148.45,0,0,92064
338,0,0,0,0,36,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),94.8,3565.65,0,20,71,19.64,2807,0,Ramona,0,0,Cable,33.044540999999995,-116.833922,0,94.8,0,0,None,33104,0,0,0,1,36,1,0.0,707.04,30.26,3565.65,1,1,92065
339,1,0,1,0,63,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,103.4,6603,1,61,14,48.95,4352,1,San Diego,1,1,Cable,32.85723,-117.209774,1,107.53600000000002,0,2,None,34902,0,0,1,1,63,3,92.44,3083.850000000001,0.0,6603.0,0,1,92122
340,0,1,0,0,32,1,0,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),54.65,1830.1,0,69,14,19.92,4045,0,Rancho Santa Fe,0,0,Cable,33.012751,-117.200617,0,54.65,0,0,None,7615,1,0,0,0,32,0,256.0,637.44,0.0,1830.1,0,0,92067
341,0,0,1,0,71,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),85.75,6223.8,0,59,18,30.68,4487,0,San Marcos,1,0,DSL,33.162624,-117.17086299999998,1,85.75,0,3,None,52664,1,0,1,1,71,1,1120.0,2178.28,4.6,6223.8,0,0,92069
342,0,0,1,1,66,1,1,DSL,1,1,0,0,Month-to-month,1,Bank transfer (automatic),67.45,4508.65,0,22,59,23.2,4172,0,Santa Ysabel,1,0,Fiber Optic,33.174725,-116.743329,1,67.45,1,6,None,1143,0,0,1,0,66,1,2660.0,1531.2,41.67,4508.65,1,0,92070
343,1,0,0,0,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.5,1328.15,0,50,0,35.35,5997,0,Santee,0,1,NA,32.847336,-116.99760500000001,0,20.5,0,0,None,53510,0,0,0,0,63,3,0.0,2227.05,15.62,1328.15,0,0,92071
344,0,0,0,1,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.25,865,0,39,0,6.61,3972,0,Solana Beach,0,0,NA,33.001813,-117.263628,0,20.25,0,0,None,12173,0,2,0,0,41,2,0.0,271.01,46.78,865.0,0,0,92075
345,0,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,72.1,72.1,0,72,22,7.77,4432,0,San Marcos,0,0,DSL,33.119028,-117.166036,0,72.1,0,0,Offer E,6760,0,0,0,0,1,3,0.0,7.77,0.0,72.1,0,1,92078
346,0,0,0,0,2,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.4,168.2,1,47,9,10.53,4157,1,San Diego,0,0,Cable,32.85723,-117.209774,0,94.016,0,0,Offer E,34902,0,0,0,1,2,4,0.0,21.06,0.0,168.2,0,1,92122
347,0,0,1,0,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.45,1303.5,0,26,0,23.52,5540,0,Vista,0,0,NA,33.17494,-117.24276100000002,1,19.45,0,9,None,62036,0,0,1,0,70,0,0.0,1646.4,14.49,1303.5,1,0,92083
348,0,0,0,0,23,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,44.95,996.85,0,47,14,0.0,3248,0,Vista,0,0,DSL,33.22784,-117.200024,0,44.95,0,0,None,44692,0,0,0,1,23,1,140.0,0.0,25.84,996.85,0,0,92084
349,0,1,1,0,64,1,0,Fiber optic,1,1,0,1,One year,0,Bank transfer (automatic),97.0,6430.9,0,69,11,3.76,4053,0,Warner Springs,1,0,Fiber Optic,33.323705,-116.626907,1,97.0,0,9,None,1205,0,0,1,0,64,0,0.0,240.64,0.0,6430.9,0,1,92086
350,1,0,1,1,37,1,1,DSL,1,0,0,0,Two year,1,Credit card (automatic),62.8,2278.75,0,57,9,4.5,5229,0,Rancho Santa Fe,1,1,DSL,32.993559999999995,-117.207121,1,62.8,0,6,None,1072,1,0,1,0,37,1,0.0,166.5,16.97,2278.75,0,1,92091
351,1,0,0,1,17,1,0,DSL,0,0,0,0,One year,0,Mailed check,44.6,681.4,0,27,73,13.02,2130,0,San Diego,0,1,DSL,32.725229999999996,-117.171346,0,44.6,0,0,None,27505,0,1,0,0,17,1,0.0,221.34,0.0,681.4,1,1,92101
352,0,1,0,0,7,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.15,574.35,0,72,28,16.36,2415,0,San Diego,0,0,Fiber Optic,32.716007,-117.11746200000002,0,89.15,0,0,None,47140,0,0,0,0,7,1,161.0,114.52,0.0,574.35,0,0,92102
353,1,0,1,1,4,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),84.8,371.9,1,26,21,28.77,4939,1,San Diego,1,1,Cable,32.85723,-117.209774,1,88.19200000000001,0,5,Offer E,34902,0,0,1,1,4,1,78.0,115.08,0.0,371.9,1,0,92122
354,0,1,0,0,21,0,No phone service,DSL,1,0,1,0,Month-to-month,1,Electronic check,41.9,840.1,1,77,9,0.0,4778,1,San Diego,0,0,DSL,32.85723,-117.209774,0,43.576,0,0,None,34902,0,0,0,0,21,2,0.0,0.0,0.0,840.1,0,1,92122
355,0,0,0,0,10,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),80.25,846,1,40,12,27.1,3598,1,San Diego,0,0,Fiber Optic,32.85723,-117.209774,0,83.46000000000002,0,0,None,34902,0,0,0,1,10,2,102.0,271.0,0.0,846.0,0,0,92122
356,0,1,0,0,16,1,1,DSL,1,0,0,0,Month-to-month,1,Electronic check,54.1,889,0,70,29,9.72,2276,0,San Diego,0,0,Fiber Optic,32.71346,-117.236378,0,54.1,0,0,Offer D,18525,0,0,0,0,16,1,0.0,155.52,0.0,889.0,0,1,92106
357,1,0,1,0,64,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,105.25,6823.4,0,29,30,40.18,5682,0,San Diego,0,1,Fiber Optic,32.741852,-117.243453,1,105.25,0,5,None,27959,1,0,1,1,64,1,204.7,2571.52,23.67,6823.4,1,1,92107
358,1,1,1,0,27,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),30.75,805.1,1,71,14,0.0,2927,1,San Diego,0,1,DSL,32.85723,-117.209774,1,31.98,0,0,None,34902,0,0,0,0,27,2,113.0,0.0,0.0,805.1,0,0,92122
359,1,0,1,1,42,1,1,Fiber optic,1,0,1,1,One year,0,Electronic check,97.1,4016.75,0,62,23,13.23,2170,0,San Diego,0,1,Fiber Optic,32.787836,-117.232376,1,97.1,0,1,None,46086,0,0,1,1,42,2,924.0,555.66,46.56,4016.75,0,0,92109
360,1,0,0,1,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.2,83.75,0,59,0,12.22,5169,0,San Diego,0,1,NA,32.76501,-117.19938,0,20.2,1,0,Offer E,24169,0,0,0,0,5,0,0.0,61.1,0.0,83.75,0,0,92110
361,0,0,0,0,41,1,0,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),98.8,3959.15,0,64,2,10.26,5584,0,San Diego,0,0,Fiber Optic,32.805518,-117.16905200000001,0,98.8,0,0,None,46828,1,0,0,1,41,0,0.0,420.66,27.09,3959.15,0,1,92111
362,1,0,1,0,58,1,0,DSL,0,0,0,0,One year,0,Credit card (automatic),50.3,2878.55,0,61,18,18.37,5232,0,San Diego,1,1,Fiber Optic,32.697098,-117.11658700000001,1,50.3,0,10,None,47431,0,0,1,0,58,3,0.0,1065.46,10.23,2878.55,0,1,92113
363,0,0,0,0,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.55,945.7,0,34,0,44.69,5404,0,San Diego,0,0,NA,32.707892,-117.05512,0,20.55,0,0,None,66838,0,1,0,0,47,2,0.0,2100.43,0.0,945.7,0,0,92114
364,1,0,0,0,18,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.9,1373.05,0,51,20,26.84,4668,0,San Diego,0,1,Fiber Optic,32.762506,-117.07245,0,75.9,0,0,None,56887,1,0,0,0,18,0,275.0,483.12,15.57,1373.05,0,0,92115
365,1,0,0,0,5,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),96.5,492.55,1,54,9,20.86,5383,1,San Diego,1,1,Cable,32.85723,-117.209774,0,100.36,0,0,Offer E,34902,0,0,0,1,5,4,44.0,104.3,0.0,492.55,0,0,92122
366,1,0,1,0,23,1,0,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),59.95,1406,0,25,69,3.67,5379,0,San Diego,0,1,DSL,32.825086,-117.199424,1,59.95,0,5,None,51213,0,0,1,1,23,1,970.0,84.41,26.55,1406.0,1,0,92117
367,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.15,19.15,0,35,0,22.37,2577,0,Coronado,0,0,NA,32.68674,-117.18661200000001,0,19.15,0,0,None,24093,0,0,0,0,1,0,0.0,22.37,0.0,19.15,0,0,92118
368,1,0,1,0,71,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),98.65,6962.85,0,60,10,34.72,5101,0,San Diego,1,1,DSL,32.802959,-117.02709499999999,1,98.65,0,8,None,21866,0,0,1,1,71,0,696.0,2465.12,0.0,6962.85,0,0,92119
369,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),112.6,8126.65,0,47,14,17.3,6486,0,San Diego,1,1,Fiber Optic,32.807867,-117.060993,1,112.6,1,2,None,25569,1,0,1,1,72,3,0.0,1245.6,0.0,8126.65,0,1,92120
370,1,0,1,1,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.6,690.25,0,63,0,34.22,5212,0,San Diego,0,1,NA,32.898613,-117.202937,1,20.6,0,2,None,4258,0,0,1,0,33,0,0.0,1129.26,0.0,690.25,0,0,92121
371,1,0,0,0,2,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.65,181.5,1,22,30,40.43,3878,1,San Diego,0,1,Fiber Optic,32.85723,-117.209774,0,89.07600000000002,0,0,Offer E,34902,0,0,0,1,2,0,54.0,80.86,0.0,181.5,1,0,92122
372,1,0,0,1,24,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,35.75,830.8,0,44,20,0.0,5531,0,San Diego,0,1,Fiber Optic,32.808814,-117.134694,0,35.75,0,0,None,25232,1,0,0,0,24,2,0.0,0.0,0.0,830.8,0,1,92123
373,0,0,1,1,56,1,1,Fiber optic,0,1,0,1,One year,1,Credit card (automatic),99.75,5608.4,0,45,19,20.53,5926,0,San Diego,1,0,DSL,32.827238,-117.08928700000001,1,99.75,0,9,None,30206,1,0,1,1,56,2,0.0,1149.68,0.0,5608.4,0,1,92124
374,1,0,0,0,37,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),96.1,3646.8,0,28,41,21.84,2640,0,San Diego,0,1,DSL,32.886925,-117.152162,0,96.1,0,0,None,74232,0,0,0,1,37,0,0.0,808.08,0.0,3646.8,1,1,92126
375,0,0,0,0,43,1,1,DSL,0,1,1,1,One year,0,Credit card (automatic),85.1,3662.25,0,29,53,2.49,2319,0,San Diego,1,0,Fiber Optic,33.017518,-117.11845600000001,0,85.1,0,0,None,20046,1,0,0,1,43,0,1941.0,107.07,0.0,3662.25,1,0,92127
376,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,25.35,25.35,0,31,13,0.0,4193,0,San Diego,0,1,Fiber Optic,33.000269,-117.072093,0,25.35,0,0,None,42733,0,0,0,0,1,1,0.0,0.0,0.0,25.35,0,1,92128
377,0,0,1,0,25,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),104.95,2566.5,1,48,11,8.91,3642,1,San Diego,1,0,Cable,32.85723,-117.209774,1,109.148,0,1,Offer C,34902,1,1,1,1,25,3,0.0,222.75,0.0,2566.5,0,1,92122
378,0,0,0,0,61,1,1,DSL,1,1,1,1,Two year,0,Electronic check,89.65,5308.7,0,52,8,23.45,6149,0,San Diego,1,0,DSL,32.957195,-117.202542,0,89.65,0,0,None,28201,1,0,0,1,61,1,425.0,1430.45,0.0,5308.7,0,0,92130
379,1,0,0,0,17,1,1,Fiber optic,0,0,0,0,One year,0,Electronic check,86.75,1410.25,0,41,4,49.71,5863,0,San Diego,1,1,Fiber Optic,32.89325,-117.08709099999999,0,86.75,0,0,None,29283,1,0,0,0,17,1,56.0,845.07,0.0,1410.25,0,0,92131
380,0,0,1,0,41,1,0,Fiber optic,0,1,0,0,One year,1,Bank transfer (automatic),86.2,3339.05,0,53,16,13.23,5325,0,San Diego,1,0,Cable,32.677716,-117.04766599999999,1,86.2,0,3,None,36351,1,0,1,0,41,0,0.0,542.4300000000002,0.0,3339.05,0,1,92139
381,1,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,50.65,50.65,1,26,65,14.78,2431,1,San Diego,0,1,DSL,32.85723,-117.209774,0,52.676,0,0,Offer E,34902,0,1,0,1,1,1,0.0,14.78,0.0,50.65,1,0,92122
382,1,1,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),64.8,4732.35,0,78,24,0.0,4886,0,San Ysidro,1,1,DSL,32.555828000000005,-117.04007299999999,1,64.8,0,1,Offer A,28488,1,0,1,0,72,1,0.0,0.0,0.0,4732.35,0,1,92173
383,1,0,0,0,1,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),90.85,90.85,1,64,26,8.56,3424,1,San Diego,0,1,DSL,32.85723,-117.209774,0,94.484,0,0,Offer E,34902,0,0,0,1,1,2,0.0,8.56,0.0,90.85,0,1,92122
384,1,0,0,0,48,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),108.1,5067.45,0,59,4,9.91,5994,0,Indio,1,1,DSL,33.752938,-116.23005500000001,0,108.1,0,0,None,2743,0,0,0,1,48,2,203.0,475.68,0.0,5067.45,0,0,92203
385,1,1,1,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,214.75,1,79,0,29.54,5888,1,San Diego,0,1,NA,32.85723,-117.209774,1,19.95,0,1,None,34902,0,0,1,0,11,2,0.0,324.94,0.0,214.75,0,0,92122
386,0,1,1,0,55,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,85.45,4874.7,1,66,30,42.82,5502,1,San Diego,1,0,DSL,32.85723,-117.209774,1,88.86800000000002,0,2,Offer B,34902,0,0,1,0,55,4,0.0,2355.1,0.0,4874.7,0,1,92122
387,0,0,0,0,42,0,No phone service,DSL,1,1,0,1,One year,1,Electronic check,54.75,2348.45,0,51,13,0.0,3179,0,Banning,1,0,Fiber Optic,33.936298,-116.849577,0,54.75,0,0,None,25859,1,0,0,1,42,0,0.0,0.0,0.0,2348.45,0,1,92220
388,1,0,0,0,44,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Mailed check,90.4,4063,0,50,16,44.92,4751,0,Beaumont,1,1,Fiber Optic,33.946982,-116.977672,0,90.4,0,0,None,17721,0,0,0,1,44,1,0.0,1976.48,0.0,4063.0,0,1,92223
389,1,0,0,1,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.0,44,0,62,29,15.66,4020,0,Blythe,0,1,Fiber Optic,33.674583,-114.71611999999999,0,44.0,2,0,None,24659,0,0,0,0,1,0,0.0,15.66,0.0,44.0,0,0,92225
390,0,0,0,0,27,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.6,2595.25,0,49,24,35.17,2026,0,Brawley,0,0,Fiber Optic,33.03933,-115.19185700000001,0,95.6,0,0,None,23394,0,0,0,1,27,0,62.29,949.59,0.0,2595.25,0,1,92227
391,1,1,1,0,27,1,1,DSL,0,1,1,1,Month-to-month,1,Bank transfer (automatic),84.8,2309.55,0,77,21,33.57,5352,0,Cabazon,1,1,Cable,33.929812,-116.76058,1,84.8,0,5,None,2355,1,0,1,0,27,0,48.5,906.39,0.0,2309.55,0,1,92230
392,0,1,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.3,89.3,0,73,22,23.91,3805,0,Calexico,0,0,DSL,32.690653999999995,-115.431225,0,44.3,0,0,Offer E,27804,0,0,0,0,2,0,20.0,47.82,0.0,89.3,0,0,92231
393,0,0,0,0,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,367.55,0,47,0,32.03,3245,0,Calipatria,0,0,NA,33.143826000000004,-115.49748500000001,0,19.9,0,0,None,7857,0,0,0,0,19,2,0.0,608.57,0.0,367.55,0,0,92233
394,0,1,1,0,42,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.05,3944.5,0,76,10,42.29,2677,0,Cathedral City,0,0,Fiber Optic,33.829583,-116.474131,1,95.05,0,10,None,43141,0,0,1,0,42,2,0.0,1776.18,0.0,3944.5,0,1,92234
395,0,0,0,0,66,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),90.05,5965.95,0,61,24,13.28,5813,0,Coachella,1,0,Fiber Optic,33.680031,-116.171678,0,90.05,0,0,None,23170,1,0,0,1,66,0,1432.0,876.4799999999998,0.0,5965.95,0,0,92236
396,1,1,1,0,33,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),109.9,3694.7,0,78,20,25.15,5655,0,Desert Center,1,1,Fiber Optic,33.889604999999996,-115.25700900000001,1,109.9,0,7,None,964,1,0,1,0,33,0,0.0,829.9499999999998,0.0,3694.7,0,1,92239
397,0,0,0,0,34,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),73.95,2524.45,1,63,15,1.55,5795,1,San Diego,0,0,Fiber Optic,32.85723,-117.209774,0,76.908,0,0,Offer C,34902,0,0,0,0,34,0,379.0,52.7,0.0,2524.45,0,0,92122
398,1,1,0,0,33,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,54.6,1803.7,0,74,11,0.0,5322,0,Desert Hot Springs,1,1,Fiber Optic,33.832799,-116.250973,0,54.6,0,0,Offer C,5529,1,0,0,0,33,0,198.0,0.0,0.0,1803.7,0,0,92241
399,0,0,1,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.05,415.1,0,44,0,17.82,3742,0,Earp,0,0,NA,34.137741999999996,-114.36514,1,20.05,0,10,None,1564,0,1,1,0,23,1,0.0,409.86,0.0,415.1,0,0,92242
400,0,0,0,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.75,624.15,0,46,0,43.8,4691,0,El Centro,0,0,NA,32.770393,-115.60915,0,19.75,0,0,None,43712,0,0,0,0,32,0,0.0,1401.6,0.0,624.15,0,0,92243
401,0,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.05,237.7,0,52,0,26.85,5355,0,Heber,0,0,NA,32.730583,-115.50108300000001,0,20.05,0,0,None,3535,0,0,0,0,11,4,0.0,295.35,0.0,237.7,0,0,92249
402,1,0,1,1,69,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),99.45,7007.6,1,30,29,48.8,4020,1,San Diego,1,1,DSL,32.85723,-117.209774,1,103.428,0,2,Offer A,34902,0,0,1,1,69,2,2032.0,3367.2,0.0,7007.6,0,0,92122
403,0,0,1,0,68,1,0,DSL,1,0,0,0,One year,0,Bank transfer (automatic),55.9,3848.8,0,49,14,44.79,5160,0,Imperial,0,0,Cable,32.858595,-115.662709,1,55.9,0,9,None,14546,1,0,1,0,68,1,539.0,3045.72,0.0,3848.8,0,0,92251
404,1,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.7,419.4,0,62,0,27.11,2120,0,Joshua Tree,0,1,NA,34.167235999999995,-116.28151100000001,0,19.7,0,0,None,8141,0,0,0,0,20,1,0.0,542.2,0.0,419.4,0,0,92252
405,1,0,0,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.8,1468.75,0,39,0,30.44,5368,0,La Quinta,0,1,NA,33.695532,-116.310571,0,19.8,0,0,Offer A,23971,0,0,0,0,72,1,0.0,2191.6800000000007,0.0,1468.75,0,0,92253
406,1,0,1,1,60,1,1,Fiber optic,1,0,1,0,One year,1,Bank transfer (automatic),95.4,5812,0,59,29,5.43,4149,0,Mecca,1,1,DSL,33.543834999999994,-115.99390600000001,1,95.4,0,5,Offer B,8768,0,1,1,0,60,2,0.0,325.7999999999999,0.0,5812.0,0,1,92254
407,1,1,1,1,32,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Mailed check,93.95,2861.45,0,71,23,31.86,2844,0,Morongo Valley,0,1,Fiber Optic,34.097863000000004,-116.59456100000001,1,93.95,1,9,Offer C,3499,0,0,1,1,32,2,658.0,1019.52,0.0,2861.45,0,0,92256
408,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.9,19.9,1,59,0,36.63,3351,1,San Diego,0,0,NA,32.85723,-117.209774,0,19.9,0,0,Offer E,34902,0,0,0,0,1,2,0.0,36.63,0.0,19.9,0,0,92122
409,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.6,19.6,1,52,0,14.17,3448,1,San Diego,0,1,NA,32.85723,-117.209774,0,19.6,0,0,Offer E,34902,0,0,0,0,1,5,0.0,14.17,0.0,19.6,0,0,92122
410,1,1,0,0,3,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,81.35,233.7,1,77,15,9.22,2818,1,San Diego,0,1,Cable,32.85723,-117.209774,0,84.604,0,0,Offer E,34902,0,3,0,0,3,1,3.51,27.660000000000004,0.0,233.7,0,1,92122
411,0,0,1,0,46,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),24.45,1066.15,0,55,0,35.46,2438,0,Palm Desert,0,0,NA,33.694501,-116.41271100000002,1,24.45,0,9,Offer B,29340,0,0,1,0,46,1,0.0,1631.16,0.0,1066.15,0,0,92260
412,0,0,1,0,29,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.95,2149.05,0,62,17,5.39,3483,0,Palm Springs,0,0,Cable,33.839989,-116.65921499999999,1,74.95,0,3,None,24924,0,0,1,0,29,2,0.0,156.31,0.0,2149.05,0,1,92262
413,1,0,0,0,51,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,87.35,4473,0,21,52,1.51,4899,0,Palm Springs,1,1,DSL,33.745746000000004,-116.514215,0,87.35,0,0,Offer B,18884,1,1,0,0,51,2,0.0,77.01,0.0,4473.0,1,1,92264
414,0,1,1,0,48,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),70.65,3545.05,0,72,21,12.6,5523,0,Palo Verde,0,0,DSL,33.3249,-114.758334,1,70.65,0,10,None,291,0,0,1,0,48,2,0.0,604.8,0.0,3545.05,0,1,92266
415,0,0,1,1,16,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),73.25,1195.75,0,58,20,40.03,3624,0,Parker Dam,0,0,Fiber Optic,34.273872,-114.192901,1,73.25,1,6,Offer D,131,0,0,1,0,16,1,239.0,640.48,0.0,1195.75,0,0,92267
416,1,0,1,0,70,1,1,Fiber optic,0,1,0,1,Two year,1,Bank transfer (automatic),98.7,6858.9,0,23,42,45.24,5582,0,Pioneertown,1,1,Cable,34.201108000000005,-116.593456,1,98.7,0,5,Offer A,354,1,2,1,1,70,1,0.0,3166.8,0.0,6858.9,1,1,92268
417,0,0,1,1,40,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.8,1024.7,0,27,0,33.44,3021,0,Rancho Mirage,0,0,NA,33.763678000000006,-116.429928,1,24.8,2,2,Offer B,12465,0,1,1,0,40,1,0.0,1337.6,0.0,1024.7,1,0,92270
418,0,0,1,1,22,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,83.3,1845.9,1,23,58,4.01,3804,1,Seeley,0,0,Cable,32.790282,-115.689559,1,86.632,0,4,None,1632,0,0,1,1,22,0,1071.0,88.22,0.0,1845.9,1,0,92273
419,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.3,75.3,1,80,19,35.09,4902,1,Thermal,1,0,Cable,33.53604,-116.119222,0,78.312,0,0,Offer E,17018,0,1,0,0,1,7,0.0,35.09,0.0,75.3,0,1,92274
420,0,0,1,1,5,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,24.3,132.25,0,41,0,6.7,3181,0,Salton City,0,0,NA,33.28156,-115.955541,1,24.3,3,6,None,799,0,0,1,0,5,1,0.0,33.5,0.0,132.25,0,0,92275
421,0,0,0,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.85,515.45,0,61,4,27.46,5501,0,Thousand Palms,0,0,Fiber Optic,33.849263,-116.382778,0,69.85,0,0,None,6242,0,0,0,0,7,1,21.0,192.22,0.0,515.45,0,0,92276
422,1,0,0,1,29,1,1,Fiber optic,0,1,0,1,One year,0,Credit card (automatic),100.55,2830.45,0,46,23,49.92,3055,0,Escondido,1,1,Fiber Optic,33.141265000000004,-116.967221,0,100.55,0,0,None,48690,1,0,0,1,29,0,651.0,1447.68,0.0,2830.45,0,0,92027
423,1,0,1,1,44,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,25.7,1110.5,0,54,0,15.33,3037,0,Twentynine Palms,0,1,NA,34.457829,-116.13958899999999,1,25.7,0,10,Offer B,14104,0,0,1,0,44,1,0.0,674.52,0.0,1110.5,0,0,92278
424,0,0,0,0,10,0,No phone service,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),40.7,449.3,0,31,24,0.0,2164,0,Escondido,1,0,DSL,33.141265000000004,-116.967221,0,40.7,0,0,Offer D,48690,0,0,0,0,10,2,0.0,0.0,0.0,449.3,0,1,92027
425,0,1,1,0,55,1,1,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),51.65,2838.55,0,75,29,29.53,4763,0,Westmorland,0,0,DSL,33.03679,-115.60503,1,51.65,0,5,None,2388,0,0,1,0,55,2,82.32,1624.15,0.0,2838.55,0,1,92281
426,1,1,1,0,52,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),105.1,5376.4,0,79,9,29.15,4621,0,White Water,1,1,Fiber Optic,33.972293,-116.654195,1,105.1,0,4,None,805,0,0,1,1,52,0,484.0,1515.8,0.0,5376.4,0,0,92282
427,0,0,1,1,10,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,85.95,858.6,0,20,76,6.5,4922,0,Winterhaven,0,0,Cable,32.852947,-114.850784,1,85.95,2,0,Offer D,3663,0,0,0,1,10,0,653.0,65.0,0.0,858.6,1,0,92283
428,1,0,0,0,18,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.6,1395.05,0,27,42,15.18,4030,0,Yucca Valley,0,1,Fiber Optic,34.159534,-116.42598400000001,0,75.6,0,0,Offer D,20486,0,1,0,0,18,1,0.0,273.24,0.0,1395.05,1,1,92284
429,0,0,1,0,68,1,1,DSL,1,0,0,0,One year,0,Bank transfer (automatic),58.25,3975.7,0,49,30,41.46,4620,0,Landers,0,0,Cable,34.341737,-116.53941599999999,1,58.25,0,4,Offer A,2182,1,2,1,0,68,4,1193.0,2819.28,0.0,3975.7,0,0,92285
430,0,0,1,1,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.4,1182.55,1,22,0,46.27,4221,1,Adelanto,0,0,NA,34.667815000000004,-117.53618300000001,1,19.4,0,3,None,18980,0,0,1,0,61,4,0.0,2822.4700000000007,0.0,1182.55,1,0,92301
431,0,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,1,Credit card (automatic),65.2,4784.45,0,56,30,0.0,5092,0,Amboy,1,0,DSL,34.559882,-115.63716399999998,1,65.2,0,5,Offer A,42,1,0,1,1,72,1,143.53,0.0,0.0,4784.45,0,1,92304
432,1,0,0,0,2,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,53.45,119.5,0,30,76,12.59,3477,0,Angelus Oaks,1,1,Fiber Optic,34.1678,-116.86433000000001,0,53.45,0,0,None,301,0,0,0,0,2,2,91.0,25.18,0.0,119.5,0,0,92305
433,1,0,0,0,12,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),45.4,518.9,1,49,15,11.12,2887,1,Fallbrook,0,1,DSL,33.362575,-117.299644,0,47.216,0,0,None,42239,0,0,0,0,12,4,78.0,133.44,0.0,518.9,0,0,92028
434,1,0,1,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Electronic check,19.75,899.45,0,21,0,35.46,2011,0,Apple Valley,0,1,NA,34.424926,-117.184503,1,19.75,0,1,Offer B,28819,0,1,1,0,41,1,0.0,1453.86,0.0,899.45,1,0,92308
435,0,0,0,0,26,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),44.45,1183.8,0,46,29,0.0,3080,0,Baker,1,0,DSL,35.28952,-116.09221399999998,0,44.45,0,0,None,904,1,0,0,0,26,1,343.0,0.0,0.0,1183.8,0,0,92309
436,1,0,1,0,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.85,720.05,0,26,0,12.61,5744,0,Fort Irwin,0,1,NA,35.349241,-116.77028100000001,1,20.85,0,1,None,9465,0,1,1,0,36,2,0.0,453.96,0.0,720.05,1,0,92310
437,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),114.05,8468.2,0,52,3,30.75,4842,0,Barstow,1,1,Fiber Optic,34.965648,-117.00150900000001,1,114.05,0,5,Offer A,31293,1,0,1,1,72,0,254.0,2214.0,0.0,8468.2,0,0,92311
438,1,0,1,0,35,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),89.85,3161.2,0,30,51,24.83,4945,0,Grand Terrace,0,1,Fiber Optic,34.029175,-117.30721100000001,1,89.85,0,0,None,11024,1,0,0,1,35,2,0.0,869.05,0.0,3161.2,0,1,92313
439,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,55.05,55.05,0,59,15,14.65,2962,0,Big Bear City,1,1,DSL,34.278967,-116.773825,0,55.05,0,0,None,9899,1,0,0,0,1,1,0.0,14.65,0.0,55.05,0,1,92314
440,0,0,1,1,16,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,112.95,1882.55,0,49,12,46.45,2683,0,Big Bear Lake,1,0,Fiber Optic,34.242058,-116.89801999999999,1,112.95,1,8,Offer D,5447,1,0,1,1,16,1,0.0,743.2,0.0,1882.55,0,1,92315
441,0,1,0,0,49,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Credit card (automatic),101.55,5070.4,0,76,14,24.84,5348,0,Bloomington,0,0,Fiber Optic,34.059722,-117.39103999999999,0,101.55,0,0,None,25995,0,0,0,1,49,2,0.0,1217.16,0.0,5070.4,0,1,92316
442,0,0,1,0,54,1,1,Fiber optic,1,1,1,1,One year,1,Mailed check,114.65,6049.5,0,63,26,11.4,4488,0,Calimesa,1,0,Fiber Optic,33.982787,-117.057627,1,114.65,0,7,Offer B,7334,1,0,1,1,54,2,1573.0,615.6,0.0,6049.5,0,0,92320
443,0,0,0,1,18,1,1,DSL,1,0,0,1,Month-to-month,0,Electronic check,64.8,1166.7,0,45,28,42.45,2466,0,Cedar Glen,0,0,Fiber Optic,34.255203,-117.17565400000001,0,64.8,3,0,Offer D,455,0,0,0,1,18,1,327.0,764.1,0.0,1166.7,0,0,92321
444,0,0,1,0,36,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,80.4,2937.65,0,59,23,49.33,5544,0,Colton,0,0,DSL,34.030915,-117.273201,1,80.4,0,8,None,52202,0,0,1,1,36,0,0.0,1775.88,0.0,2937.65,0,1,92324
445,0,0,0,0,60,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.9,6396.45,1,20,78,10.7,4105,1,Crestline,1,0,DSL,34.248061,-117.29028000000001,0,110.136,0,0,None,10484,0,0,0,1,60,1,4989.0,642.0,0.0,6396.45,1,0,92325
446,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,69.55,69.55,1,54,14,29.78,2792,1,Daggett,0,0,Cable,34.875144,-116.821698,0,72.332,0,0,Offer E,678,0,2,0,0,1,3,0.0,29.78,0.0,69.55,0,0,92327
447,0,0,1,1,52,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.05,1270.25,0,30,0,5.32,5674,0,Death Valley,0,0,NA,36.27688,-117.033326,1,25.05,0,10,Offer B,443,0,0,1,0,52,1,0.0,276.64,0.0,1270.25,0,0,92328
448,1,0,1,1,8,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.75,759.55,0,26,82,22.14,5505,0,Essex,1,1,Fiber Optic,34.9436,-115.287901,1,94.75,3,4,None,115,0,1,1,1,8,1,623.0,177.12,0.0,759.55,1,0,92332
449,1,0,1,1,72,1,0,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),105.5,7611.55,0,47,19,27.25,5534,0,Fawnskin,0,1,Fiber Optic,34.274846000000004,-116.93758100000001,1,105.5,0,8,Offer A,414,1,0,1,1,72,1,0.0,1962.0,0.0,7611.55,0,1,92333
450,0,0,0,0,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,24.7,1642.75,0,53,0,4.03,5655,0,Fontana,0,0,NA,34.087558,-117.464096,0,24.7,0,0,Offer B,82630,0,0,0,0,64,0,0.0,257.92,0.0,1642.75,0,0,92335
451,0,1,0,0,22,1,0,DSL,1,0,0,1,Month-to-month,1,Mailed check,69.75,1545.4,0,78,28,49.98,3509,0,Fontana,1,0,DSL,34.136367,-117.460803,0,69.75,0,0,Offer D,54586,1,0,0,1,22,0,0.0,1099.56,0.0,1545.4,0,1,92336
452,1,0,1,0,60,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Bank transfer (automatic),60.2,3582.4,0,34,2,0.0,5359,0,Fontana,1,1,DSL,34.049671000000004,-117.468896,1,60.2,0,10,Offer B,29847,1,0,1,1,60,0,72.0,0.0,0.0,3582.4,0,0,92337
453,0,0,1,1,28,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,81.05,2227.1,1,58,14,16.85,5201,1,Ludlow,0,0,Fiber Optic,34.702766,-116.093376,1,84.292,0,1,Offer C,23,0,0,1,1,28,0,0.0,471.80000000000007,0.0,2227.1,0,1,92338
454,0,0,1,0,61,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.4,1417.9,0,20,0,20.09,4900,0,Forest Falls,0,0,NA,34.067699,-116.90389099999999,1,24.4,0,10,Offer B,958,0,0,1,0,61,0,0.0,1225.49,0.0,1417.9,1,0,92339
455,0,0,0,0,24,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.15,2494.65,0,48,4,38.79,5813,0,Green Valley Lake,1,0,Fiber Optic,34.244411,-117.072654,0,104.15,0,0,None,317,0,0,0,1,24,3,0.0,930.96,0.0,2494.65,0,1,92341
456,1,0,1,1,28,1,0,Fiber optic,0,1,1,0,One year,0,Bank transfer (automatic),92.9,2768.35,0,35,16,27.34,2037,0,Helendale,1,1,DSL,34.757783,-117.33997,1,92.9,0,1,None,4948,1,0,1,0,28,1,443.0,765.52,0.0,2768.35,0,0,92342
457,0,0,1,1,30,1,0,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),80.8,2369.3,0,24,53,15.94,4274,0,Hesperia,1,0,Cable,34.361387,-117.33750900000001,1,80.8,0,4,Offer C,68515,1,0,1,1,30,0,125.57,478.2,0.0,2369.3,1,1,92345
458,1,0,1,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,38,0,45,0,34.38,4823,0,Highland,0,1,NA,34.129677,-117.15427700000001,1,20.0,0,10,None,48245,0,0,1,0,2,2,0.0,68.76,0.0,38.0,0,0,92346
459,1,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.1,75.1,0,61,28,4.53,4120,0,Hinkley,0,1,DSL,34.983808,-117.239306,0,75.1,0,0,None,1933,0,0,0,0,1,2,0.0,4.53,0.0,75.1,0,1,92347
460,1,0,0,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,100.9,0,52,0,15.5,2231,0,Lake Arrowhead,0,1,NA,34.2565,-117.19335,0,19.65,2,0,None,9793,0,0,0,0,6,0,0.0,93.0,0.0,100.9,0,0,92352
461,0,0,1,0,24,1,0,DSL,0,1,1,1,Month-to-month,1,Bank transfer (automatic),69.45,1614.05,0,23,59,44.06,4208,0,Loma Linda,0,0,Cable,34.049315,-117.255974,1,69.45,0,8,Offer C,18068,0,0,1,1,24,0,952.0,1057.44,0.0,1614.05,1,0,92354
462,1,0,1,1,4,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,101.15,385.9,1,21,53,9.56,4417,1,Lucerne Valley,1,1,Cable,34.508417,-116.856103,1,105.196,0,3,Offer E,5256,0,1,1,1,4,3,205.0,38.24,0.0,385.9,1,0,92356
463,1,0,0,0,7,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.8,673.25,1,61,2,47.03,2031,1,Lytle Creek,0,1,Fiber Optic,34.238162,-117.534306,0,103.792,0,0,None,1090,0,2,0,1,7,3,0.0,329.2100000000001,0.0,673.25,0,1,92358
464,1,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),116.05,8404.9,0,75,13,21.37,4404,0,Mentone,1,1,DSL,34.103578000000006,-117.04054,1,116.05,0,5,Offer A,7324,1,1,1,1,72,3,0.0,1538.64,0.0,8404.9,0,1,92359
465,1,0,0,0,70,0,No phone service,DSL,0,0,0,1,Two year,1,Mailed check,40.05,2799.75,0,25,59,0.0,5055,0,Needles,0,1,Fiber Optic,34.711224,-114.702256,0,40.05,0,0,Offer A,5488,1,0,0,1,70,1,0.0,0.0,0.0,2799.75,1,1,92363
466,1,1,1,0,64,1,1,Fiber optic,0,0,1,1,Two year,0,Electronic check,102.1,6538.45,0,66,8,20.19,6270,0,Nipton,1,1,Fiber Optic,35.478736,-115.51698400000001,1,102.1,0,2,None,162,1,0,1,1,64,0,523.0,1292.16,0.0,6538.45,0,0,92364
467,1,0,1,1,72,1,1,Fiber optic,0,1,1,0,One year,1,Electronic check,89.7,6588.95,0,32,18,11.57,6016,0,Temecula,0,1,Cable,33.507255,-117.029473,1,89.7,0,2,Offer A,46171,0,2,1,0,72,2,1186.0,833.04,0.0,6588.95,0,0,92592
468,0,0,0,1,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.9,868.1,0,42,0,13.45,2809,0,Oro Grande,0,0,NA,34.647959,-117.296957,0,19.9,0,0,Offer B,909,0,0,0,0,44,0,0.0,591.8,0.0,868.1,0,0,92368
469,0,0,1,1,13,1,0,DSL,0,0,0,1,Month-to-month,0,Electronic check,55.95,734.35,1,60,30,19.05,4498,1,Phelan,0,0,Cable,34.441123,-117.53788600000001,1,58.188,0,3,Offer D,12463,0,0,1,1,13,0,220.0,247.65,0.0,734.35,0,0,92371
470,0,1,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.65,330.6,0,71,0,24.15,4086,0,Pinon Hills,0,0,NA,34.459322,-117.629729,0,20.65,0,0,Offer D,4280,0,0,0,0,17,1,0.0,410.55,0.0,330.6,0,0,92372
471,1,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.0,55,1,25,58,47.22,4877,1,Redlands,0,1,Cable,34.003243,-117.13828600000001,0,57.2,0,0,None,31230,0,2,0,1,1,3,0.0,47.22,0.0,55.0,1,0,92373
472,1,0,1,0,9,1,0,DSL,0,0,1,1,Month-to-month,1,Mailed check,70.05,564.4,0,24,82,14.91,4900,0,Redlands,1,1,DSL,34.064073,-117.16615800000001,1,70.05,0,2,None,36675,0,0,1,1,9,0,463.0,134.19,0.0,564.4,1,0,92374
473,1,0,1,0,24,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,53.6,1315.35,0,56,3,1.02,2977,0,Rialto,0,1,DSL,34.109775,-117.378904,1,53.6,0,7,Offer C,75882,1,0,1,0,24,1,0.0,24.48,0.0,1315.35,0,1,92376
474,0,0,1,1,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.7,74.7,1,52,9,21.91,5980,1,Rialto,0,0,Cable,34.156758,-117.40468600000001,1,77.688,0,0,None,18518,0,1,0,0,1,4,0.0,21.91,0.0,74.7,0,0,92377
475,1,0,0,0,24,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.25,1861.5,1,52,22,49.3,4418,1,Running Springs,0,1,Cable,34.186211,-117.07683,0,83.46000000000002,0,0,Offer C,5395,0,5,0,0,24,1,410.0,1183.1999999999996,0.0,1861.5,0,0,92382
476,1,1,1,1,35,1,0,DSL,0,1,1,1,Month-to-month,1,Electronic check,76.05,2747.2,0,77,17,14.19,5479,0,Shoshone,0,1,Fiber Optic,35.924252,-116.18866799999999,1,76.05,1,6,Offer C,87,1,0,1,1,35,0,0.0,496.65,0.0,2747.2,0,1,92384
477,0,0,1,1,7,1,0,DSL,1,1,1,0,Month-to-month,1,Electronic check,75.7,554.05,0,47,53,16.22,2950,0,Sugarloaf,1,0,Cable,34.243088,-116.83001499999999,1,75.7,3,8,None,1834,1,0,1,0,7,3,294.0,113.54,0.0,554.05,0,0,92386
478,1,0,0,0,5,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.1,453.4,1,61,12,31.09,4192,1,Fallbrook,0,1,Cable,33.362575,-117.299644,0,99.944,0,0,None,42239,1,0,0,1,5,7,54.0,155.45,0.0,453.4,0,0,92028
479,0,0,0,1,15,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),69.0,994.8,1,40,31,4.67,5671,1,Victorville,0,0,DSL,34.486835,-117.362274,0,71.76,0,0,Offer D,63235,0,2,0,0,15,6,0.0,70.05,0.0,994.8,0,1,92392
480,1,0,1,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.65,225.75,0,48,0,40.76,3372,0,Victorville,0,1,NA,34.567058,-117.362329,1,19.65,2,2,Offer D,12083,0,0,1,0,11,1,0.0,448.36,0.0,225.75,0,0,92394
481,0,0,1,0,48,0,No phone service,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),45.3,2145,1,28,64,0.0,4926,1,Wrightwood,1,0,Cable,34.358321000000004,-117.61826299999998,1,47.111999999999995,0,3,None,4253,0,0,1,1,48,3,0.0,0.0,0.0,2145.0,1,1,92397
482,0,1,0,0,20,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,81.45,1671.6,0,74,21,23.18,2416,0,Yermo,0,0,Fiber Optic,35.013298999999996,-116.834092,0,81.45,0,0,Offer D,1195,0,0,0,1,20,1,351.0,463.6,0.0,1671.6,0,0,92398
483,0,0,1,0,72,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),108.5,8003.8,0,50,16,38.44,6288,0,Yucaipa,1,0,Fiber Optic,34.045970000000004,-117.011825,1,108.5,0,2,Offer A,41575,1,0,1,1,72,2,1281.0,2767.68,0.0,8003.8,0,0,92399
484,0,0,1,1,8,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,83.55,680.05,1,32,28,32.32,2879,1,San Bernardino,0,0,Cable,34.105934999999995,-117.2914,1,86.89200000000001,0,1,None,1779,0,1,1,0,8,2,190.0,258.56,0.0,680.05,0,0,92401
485,1,0,1,1,72,1,1,Fiber optic,0,0,0,1,Two year,1,Credit card (automatic),84.5,6130.85,0,62,20,44.0,6202,0,San Bernardino,0,1,Cable,34.183285999999995,-117.221722,1,84.5,2,4,Offer A,53636,0,0,1,1,72,1,122.62,3168.0,0.0,6130.85,0,1,92404
486,0,0,0,0,15,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.15,1415,0,64,28,32.07,2565,0,San Bernardino,0,0,Cable,34.142747,-117.30086399999999,0,100.15,0,0,Offer D,24644,0,0,0,1,15,0,0.0,481.05,0.0,1415.0,0,1,92405
487,1,0,0,0,72,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),88.6,6201.95,0,26,48,44.46,5842,0,San Bernardino,1,1,Cable,34.250069,-117.39394899999999,0,88.6,0,0,Offer A,49355,1,1,0,1,72,1,0.0,3201.12,0.0,6201.95,1,1,92407
488,0,0,1,1,0,0,No phone service,DSL,1,0,1,0,Two year,1,Bank transfer (automatic),52.55, ,0,43,20,0.0,2578,0,San Bernardino,1,0,DSL,34.084909,-117.25810700000001,1,52.55,0,2,None,12149,1,0,1,0,10,0,0.0,0.0,0.0,525.5,0,1,92408
489,1,0,0,1,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.35,74.35,1,32,2,14.02,2814,1,San Bernardino,0,1,Cable,34.106922,-117.29755300000001,0,77.324,0,0,None,44556,0,2,0,0,1,3,0.0,14.02,0.0,74.35,0,0,92410
490,1,0,1,1,63,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),104.8,6597.25,0,42,76,40.73,4046,0,San Bernardino,1,1,Fiber Optic,34.122501,-117.32013799999999,1,104.8,3,4,Offer B,23146,0,1,1,1,63,1,5014.0,2565.99,0.0,6597.25,0,0,92411
491,0,0,0,0,2,1,0,DSL,0,1,1,0,Month-to-month,1,Electronic check,59.0,114.15,0,63,26,27.02,5810,0,Riverside,0,0,Fiber Optic,33.994676,-117.372498,0,59.0,0,0,None,18999,0,0,0,0,2,0,30.0,54.04,0.0,114.15,0,0,92501
492,0,0,1,0,2,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,74.4,139.4,1,28,45,9.79,4263,1,Riverside,0,0,Cable,33.890046000000005,-117.455583,1,77.376,0,1,None,71678,0,0,1,0,2,5,0.0,19.58,0.0,139.4,1,1,92503
493,1,1,1,0,61,1,1,DSL,0,1,0,1,One year,0,Bank transfer (automatic),64.05,3902.6,0,73,20,34.24,4001,0,Riverside,0,1,Fiber Optic,33.9108,-117.39815300000001,1,64.05,0,9,None,46550,0,0,1,1,61,0,781.0,2088.640000000001,0.0,3902.6,0,0,92504
494,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,20.4,0,31,0,17.81,2968,0,Riverside,0,1,NA,33.920907,-117.489426,0,20.4,0,0,None,38446,0,0,0,0,1,0,0.0,17.81,0.0,20.4,0,0,92505
495,1,0,0,0,22,0,No phone service,DSL,0,1,0,1,One year,1,Bank transfer (automatic),43.75,903.6,1,51,18,0.0,3099,1,Riverside,1,1,Cable,33.930931,-117.36178799999999,0,45.5,0,0,Offer D,42425,0,5,0,1,22,3,163.0,0.0,0.0,903.6,0,0,92506
496,1,0,1,0,28,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,60.9,1785.65,0,32,24,28.86,3851,0,Riverside,0,1,DSL,33.976328,-117.31978600000001,1,60.9,0,7,Offer C,48649,1,1,1,0,28,2,429.0,808.0799999999998,0.0,1785.65,0,0,92507
497,0,0,1,0,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.8,1397.65,0,41,0,11.71,4500,0,Riverside,0,0,NA,33.885498999999996,-117.324959,1,19.8,0,7,Offer A,17147,0,0,1,0,70,0,0.0,819.7,0.0,1397.65,0,0,92508
498,0,1,0,0,5,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,28.45,131.05,1,77,29,0.0,4099,1,Riverside,0,0,Cable,34.004379,-117.447864,0,29.588,0,0,Offer E,63999,0,0,0,0,5,4,38.0,0.0,0.0,131.05,0,0,92509
499,0,0,0,0,12,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Bank transfer (automatic),99.7,1238.45,1,49,15,16.07,2538,1,March Air Reserve Base,1,0,DSL,33.888323,-117.277533,0,103.68799999999999,0,0,Offer D,1005,0,1,0,1,12,3,186.0,192.84,0.0,1238.45,0,0,92518
500,1,0,0,0,34,1,1,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),116.25,3899.05,0,64,13,22.41,4022,0,Lake Elsinore,1,1,Cable,33.655421000000004,-117.391751,0,116.25,0,0,Offer C,38519,1,0,0,1,34,1,507.0,761.94,0.0,3899.05,0,0,92530
501,0,1,1,0,71,1,1,Fiber optic,1,0,0,0,Two year,1,Credit card (automatic),80.7,5676,0,73,17,43.99,4583,0,Lake Elsinore,0,0,Fiber Optic,33.705836,-117.31820400000001,1,80.7,0,4,Offer A,4546,0,0,1,0,71,0,96.49,3123.29,0.0,5676.0,0,1,92532
502,0,0,1,1,70,1,1,DSL,1,0,0,1,One year,0,Bank transfer (automatic),65.2,4543.15,0,50,12,29.72,6316,0,Aguanga,0,0,Fiber Optic,33.482243,-116.827173,1,65.2,0,1,Offer A,2433,0,0,1,1,70,0,545.0,2080.4,0.0,4543.15,0,0,92536
503,0,0,1,1,52,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),84.05,4326.8,0,54,26,31.96,6099,0,Anza,1,0,Cable,33.527605,-116.666551,1,84.05,2,1,Offer B,3745,1,0,1,0,52,1,0.0,1661.92,0.0,4326.8,0,1,92539
504,1,0,0,1,69,1,1,DSL,1,1,1,0,Two year,1,Credit card (automatic),79.45,5502.55,0,23,46,26.45,5189,0,Hemet,1,1,Fiber Optic,33.739415,-116.96833899999999,0,79.45,0,0,Offer A,29687,1,0,0,0,69,1,2531.0,1825.05,0.0,5502.55,1,0,92543
505,0,1,0,0,20,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,94.1,1782.4,1,77,13,48.73,2666,1,Hemet,1,0,Fiber Optic,33.644585,-116.871544,0,97.86399999999999,0,0,None,39264,0,1,0,0,20,4,232.0,974.6,0.0,1782.4,0,0,92544
506,1,0,0,1,11,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,78.0,851.8,0,63,23,47.12,4886,0,Hemet,1,1,Fiber Optic,33.734933000000005,-117.044145,0,78.0,2,0,Offer D,25694,0,0,0,0,11,1,0.0,518.3199999999998,0.0,851.8,0,1,92545
507,1,0,1,0,2,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.2,167.5,1,49,21,18.79,3715,1,Homeland,0,1,Cable,33.761894,-117.12086799999999,1,97.96799999999999,0,4,None,4283,1,0,1,1,2,2,35.0,37.58,0.0,167.5,0,0,92548
508,0,0,1,1,6,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,80.5,502.85,1,64,25,36.12,5032,1,Idyllwild,0,0,DSL,33.755039000000004,-116.741796,1,83.72,0,1,None,3588,1,2,1,0,6,4,126.0,216.72,0.0,502.85,0,0,92549
509,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,19.85,0,47,0,16.47,4905,0,Moreno Valley,0,0,NA,33.882740000000005,-117.224878,0,19.85,0,0,None,22983,0,0,0,0,1,0,0.0,16.47,0.0,19.85,0,0,92551
510,1,1,1,1,20,1,0,Fiber optic,1,0,0,1,One year,0,Credit card (automatic),94.3,1818.3,0,78,5,32.54,2574,0,Moreno Valley,1,1,Fiber Optic,33.923149,-117.244933,1,94.3,0,1,None,61205,1,0,1,0,20,1,9.09,650.8,0.0,1818.3,0,1,92553
511,1,0,0,0,61,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,106.45,6300.15,0,21,73,36.05,4842,0,Moreno Valley,1,1,DSL,33.907361,-117.109972,0,106.45,0,0,Offer B,12743,0,2,0,1,61,1,0.0,2199.05,0.0,6300.15,1,1,92555
512,0,1,1,0,5,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.35,334.8,1,72,24,45.76,5273,1,Moreno Valley,0,0,Fiber Optic,33.970661,-117.255039,1,77.324,0,4,Offer E,46214,0,2,1,0,5,4,80.0,228.8,0.0,334.8,0,0,92557
513,0,0,0,0,56,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),105.45,5916.95,0,42,3,2.5,4212,0,Mountain Center,0,0,DSL,33.638645000000004,-116.55783000000001,0,105.45,0,0,Offer B,1500,1,0,0,1,56,0,178.0,140.0,0.0,5916.95,0,0,92561
514,1,0,0,0,30,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),95.0,2852.4,0,36,29,2.87,3597,0,Murrieta,1,1,Fiber Optic,33.548869,-117.33416499999998,0,95.0,0,0,Offer C,36149,1,0,0,0,30,0,827.0,86.10000000000002,0.0,2852.4,0,0,92562
515,1,0,0,0,40,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),104.8,4131.95,1,55,9,35.58,3492,1,Murrieta,1,1,Cable,33.581045,-117.14719,0,108.992,0,0,None,18311,1,1,0,1,40,2,0.0,1423.1999999999996,0.0,4131.95,0,1,92563
516,0,0,0,0,28,1,0,DSL,1,0,0,0,One year,0,Mailed check,54.3,1546.3,0,19,48,28.42,5271,0,Nuevo,0,0,Fiber Optic,33.827690000000004,-117.102244,0,54.3,0,0,Offer C,7344,1,0,0,0,28,2,742.0,795.76,0.0,1546.3,1,0,92567
517,0,1,1,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.05,302.6,0,79,23,5.42,2064,0,Perris,0,0,Fiber Optic,33.787298,-117.320676,1,70.05,0,1,Offer E,36817,0,0,1,0,5,1,70.0,27.1,0.0,302.6,0,0,92570
518,0,1,1,0,27,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),75.2,1929.35,1,80,28,7.02,4517,1,Perris,0,0,DSL,33.828289,-117.20166599999999,1,78.20800000000001,0,2,None,26357,0,0,1,0,27,1,0.0,189.54,0.0,1929.35,0,1,92571
519,1,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.05,265.45,0,34,0,38.96,4996,0,San Jacinto,0,1,NA,33.806708,-117.02006999999999,0,20.05,0,0,Offer D,4456,0,0,0,0,12,0,0.0,467.52,0.0,265.45,0,0,92582
520,1,0,1,1,67,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,105.4,6989.45,0,37,16,38.98,5666,0,San Jacinto,1,1,Cable,33.796568,-116.924723,1,105.4,2,0,Offer A,21349,0,0,0,1,67,0,0.0,2611.66,0.0,6989.45,0,1,92583
521,1,1,1,0,29,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,51.6,1442,0,77,9,37.65,5495,0,Menifee,0,1,DSL,33.653338,-117.178271,1,51.6,0,1,Offer C,14068,0,2,1,0,29,1,12.98,1091.85,0.0,1442.0,0,1,92584
522,1,0,1,1,55,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Bank transfer (automatic),85.5,4713.4,0,29,52,41.89,6411,0,Sun City,0,1,Cable,33.739412,-117.17333400000001,1,85.5,2,1,Offer B,8692,0,0,1,1,55,0,0.0,2303.95,0.0,4713.4,1,1,92585
523,0,0,0,0,23,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),75.6,1758.6,1,47,25,27.61,2115,1,Sun City,0,0,Fiber Optic,33.707483,-117.200006,0,78.624,0,0,Offer D,18161,0,2,0,0,23,3,440.0,635.03,0.0,1758.6,0,0,92586
524,1,0,1,0,34,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.05,3480,1,22,57,23.09,2568,1,Sun City,1,1,DSL,33.69887,-117.25071000000001,1,104.052,0,2,Offer C,13151,0,0,1,1,34,5,0.0,785.06,0.0,3480.0,1,1,92587
525,1,0,0,0,52,1,0,Fiber optic,1,0,1,0,One year,0,Electronic check,91.25,4738.3,0,43,12,31.31,4770,0,Temecula,1,1,Fiber Optic,33.475493,-117.219551,0,91.25,0,0,Offer B,3070,0,0,0,0,52,0,0.0,1628.12,0.0,4738.3,0,1,92590
526,1,1,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),115.75,8399.15,0,77,17,30.78,5168,0,Temecula,1,1,Cable,33.540603999999995,-117.10909,1,115.75,1,1,Offer A,25655,1,0,1,0,72,0,142.79,2216.16,0.0,8399.15,0,1,92591
527,1,0,1,1,58,1,1,Fiber optic,0,1,1,0,One year,1,Credit card (automatic),94.7,5430.35,0,30,69,43.75,5653,0,Temecula,0,1,DSL,33.507255,-117.029473,1,94.7,3,1,Offer B,46171,1,0,1,0,58,2,3747.0,2537.5,0.0,5430.35,0,0,92592
528,1,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.6,686.95,0,52,0,20.85,3764,0,Wildomar,0,1,NA,33.617108,-117.253349,1,19.6,3,1,Offer C,19368,0,0,1,0,35,2,0.0,729.75,0.0,686.95,0,0,92595
529,0,1,0,0,56,1,1,Fiber optic,0,1,1,0,Two year,1,Bank transfer (automatic),99.9,5706.3,0,80,16,17.33,5840,0,Winchester,1,0,DSL,33.657433000000005,-117.04253999999999,0,99.9,0,0,None,4093,1,0,0,0,56,0,913.0,970.48,0.0,5706.3,0,0,92596
530,0,0,1,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),21.1,490.65,0,51,0,20.6,4368,0,Irvine,0,0,NA,33.720359,-117.733655,1,21.1,3,9,Offer C,2762,0,0,1,0,24,1,0.0,494.4,0.0,490.65,0,0,92602
531,1,0,1,1,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.05,1360.25,0,47,0,48.57,4485,0,Irvine,0,1,NA,33.688546,-117.788091,1,20.05,2,5,Offer A,27369,0,0,1,0,70,0,0.0,3399.9,0.0,1360.25,0,0,92604
532,1,0,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.95,174.45,0,25,73,37.7,5213,0,Irvine,0,1,Fiber Optic,33.703976000000004,-117.82417199999999,0,79.95,0,0,None,17621,0,0,0,0,2,1,127.0,75.4,0.0,174.45,1,0,92606
533,1,1,1,1,68,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),107.15,7379.8,0,80,12,32.11,4324,0,Foothill Ranch,1,1,DSL,33.698728,-117.67768000000001,1,107.15,1,0,Offer A,10936,1,0,0,0,68,0,0.0,2183.48,0.0,7379.8,0,1,92610
534,0,0,0,0,1,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.0,85,1,51,33,30.52,5679,1,Irvine,0,0,Fiber Optic,33.643095,-117.810896,0,88.4,0,0,Offer E,41062,0,0,0,1,1,3,0.0,30.52,0.0,85.0,0,1,92612
535,1,0,0,0,12,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,89.55,1021.75,0,60,22,33.36,2325,0,Irvine,1,1,Fiber Optic,33.680302000000005,-117.83329599999999,0,89.55,0,0,Offer D,22499,0,0,0,0,12,2,225.0,400.32,0.0,1021.75,0,0,92614
536,0,0,1,0,63,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),81.55,5029.05,0,54,24,21.15,4980,0,Irvine,0,0,Fiber Optic,33.667145,-117.73213500000001,1,81.55,0,1,Offer B,6301,0,0,1,0,63,0,1207.0,1332.4499999999996,0.0,5029.05,0,0,92618
537,0,0,1,1,33,1,0,DSL,1,1,0,0,One year,1,Mailed check,58.45,1955.4,0,24,27,8.79,4276,0,Irvine,1,0,DSL,33.716136,-117.752574,1,58.45,0,8,Offer C,26419,0,0,1,0,33,0,528.0,290.07,0.0,1955.4,1,0,92620
538,0,0,1,0,69,1,0,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),95.65,6744.2,0,32,11,46.87,5251,0,Capistrano Beach,0,0,Cable,33.458754,-117.665104,1,95.65,0,4,None,7465,0,0,1,1,69,0,742.0,3234.03,0.0,6744.2,0,0,92624
539,0,0,1,1,60,1,0,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),80.6,4946.7,0,26,42,14.0,5667,0,Corona Del Mar,1,0,Fiber Optic,33.600986999999996,-117.862734,1,80.6,0,5,None,13422,1,0,1,1,60,2,2078.0,840.0,0.0,4946.7,1,0,92625
540,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),113.1,8248.5,0,43,53,26.32,5308,0,Costa Mesa,1,0,Fiber Optic,33.678591,-117.90547099999999,1,113.1,5,10,None,48207,1,0,1,1,72,2,4372.0,1895.04,0.0,8248.5,0,0,92626
541,0,0,0,0,11,1,1,DSL,0,0,0,1,Month-to-month,1,Mailed check,58.95,601.6,0,52,10,24.57,3880,0,Costa Mesa,0,0,Cable,33.645672,-117.92261299999998,0,58.95,0,0,Offer D,62069,0,0,0,1,11,1,60.0,270.27,0.0,601.6,0,0,92627
542,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.55,19.55,0,57,0,40.63,3968,0,Dana Point,0,0,NA,33.477923,-117.70531399999999,0,19.55,0,0,None,27730,0,0,0,0,1,0,0.0,40.63,0.0,19.55,0,0,92629
543,1,0,0,0,10,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),86.05,834.1,1,33,12,5.92,2966,1,Lake Forest,0,1,DSL,33.644849,-117.68425400000001,0,89.492,0,0,Offer D,59176,0,0,0,0,10,4,100.0,59.2,0.0,834.1,0,0,92630
544,1,0,0,0,13,0,No phone service,DSL,1,0,1,0,Month-to-month,1,Credit card (automatic),45.55,597,1,52,19,0.0,4856,1,Huntington Beach,0,1,DSL,33.666301000000004,-117.969501,0,47.372,0,0,Offer D,56517,1,0,0,0,13,6,113.0,0.0,0.0,597.0,0,0,92646
545,1,0,1,1,34,1,0,Fiber optic,0,0,0,1,One year,1,Bank transfer (automatic),78.95,2647.2,0,59,12,3.54,2074,0,Huntington Beach,0,1,Fiber Optic,33.723579,-118.00544099999999,1,78.95,1,1,Offer C,58764,0,2,1,1,34,2,318.0,120.36,0.0,2647.2,0,0,92647
546,1,0,1,1,39,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Mailed check,86.3,3266,1,29,21,40.25,3364,1,Huntington Beach,0,1,Cable,33.679659,-118.016195,1,89.75200000000001,0,5,Offer C,42663,0,4,1,0,39,7,686.0,1569.75,0.0,3266.0,1,0,92648
547,0,0,0,0,65,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),105.05,6744.25,0,22,59,26.83,5742,0,Huntington Beach,0,0,DSL,33.721917,-118.043237,0,105.05,0,0,None,32304,1,0,0,1,65,0,397.91,1743.9499999999996,0.0,6744.25,1,1,92649
548,1,1,1,0,50,1,1,Fiber optic,1,1,1,0,One year,1,Bank transfer (automatic),101.9,5265.5,0,80,17,14.49,4184,0,Laguna Beach,1,1,Cable,33.570023,-117.773669,1,101.9,0,9,None,25206,0,0,1,0,50,0,895.0,724.5,0.0,5265.5,0,0,92651
549,1,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.75,311.6,0,35,0,3.49,4123,0,Laguna Hills,0,1,NA,33.606899,-117.717854,0,19.75,0,0,None,48273,0,1,0,0,15,1,0.0,52.35,0.0,311.6,0,0,92653
550,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),110.3,7966.9,0,44,51,33.01,5780,0,Midway City,1,1,Fiber Optic,33.744439,-117.98588000000001,1,110.3,4,10,None,8660,0,0,1,1,72,2,0.0,2376.72,0.0,7966.9,0,1,92655
551,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),115.6,8220.4,0,26,59,34.69,5633,0,Aliso Viejo,1,0,Fiber Optic,33.571259000000005,-117.731917,1,115.6,3,9,None,41237,1,0,1,1,72,0,4850.0,2497.68,0.0,8220.4,1,0,92656
552,1,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.35,1153.25,0,46,0,24.7,5248,0,Newport Coast,0,1,NA,33.603282,-117.82184099999999,1,19.35,2,2,None,5597,0,1,1,0,55,1,0.0,1358.5,0.0,1153.25,0,0,92657
553,0,0,1,1,23,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.6,514.75,0,27,0,25.54,5939,0,Newport Beach,0,0,NA,33.634626000000004,-117.874882,1,25.6,2,1,None,28687,0,0,1,0,23,0,0.0,587.42,0.0,514.75,1,0,92660
554,1,0,0,0,32,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.35,2596.15,1,31,23,1.49,5974,1,Newport Beach,0,1,Cable,33.601309,-117.902304,0,83.564,0,0,Offer C,4242,0,5,0,0,32,1,597.0,47.68,0.0,2596.15,0,0,92661
555,0,0,1,1,56,1,1,DSL,1,0,0,1,One year,1,Bank transfer (automatic),68.75,3808,0,58,8,42.86,6198,0,Newport Beach,1,0,Cable,33.606336,-117.893042,1,68.75,0,2,None,3124,0,0,1,1,56,0,0.0,2400.16,0.0,3808.0,0,1,92662
556,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.9,19.9,0,22,0,11.83,2010,0,Newport Beach,0,0,NA,33.62251,-117.927024,0,19.9,0,0,None,22133,0,0,0,0,1,0,0.0,11.83,0.0,19.9,1,0,92663
557,1,0,0,0,38,1,0,DSL,1,1,1,0,One year,0,Mailed check,70.6,2708.2,0,55,22,42.24,4993,0,San Clemente,0,1,Cable,33.429488,-117.60943200000001,0,70.6,0,0,Offer C,34946,1,0,0,0,38,1,0.0,1605.12,0.0,2708.2,0,1,92672
558,1,0,0,0,11,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.2,760.05,0,51,8,1.01,2535,0,San Clemente,0,1,Fiber Optic,33.4725,-117.584273,0,70.2,0,0,None,15297,0,0,0,0,11,0,61.0,11.11,0.0,760.05,0,0,92673
559,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.3,49.3,0,54,5,14.97,4209,0,San Juan Capistrano,0,1,Fiber Optic,33.521446999999995,-117.60255500000001,0,49.3,0,0,None,34321,1,0,0,0,1,0,0.0,14.97,0.0,49.3,0,1,92675
560,1,0,1,0,56,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,107.25,6033.3,0,53,25,14.43,5800,0,Silverado,0,1,Fiber Optic,33.782346000000004,-117.635263,1,107.25,0,1,None,1859,1,1,1,1,56,1,0.0,808.0799999999998,0.0,6033.3,0,1,92676
561,1,0,1,0,3,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,23.6,89.05,0,19,0,14.1,5587,0,Laguna Niguel,0,1,NA,33.529047,-117.701175,1,23.6,0,9,Offer E,62103,0,0,1,0,3,1,0.0,42.3,0.0,89.05,1,0,92677
562,1,0,1,1,7,1,0,DSL,1,0,1,1,Month-to-month,0,Credit card (automatic),69.7,516.15,0,63,51,5.17,4326,0,Trabuco Canyon,0,1,Cable,33.631119,-117.567346,1,69.7,3,6,Offer E,32268,0,0,1,1,7,1,0.0,36.19,0.0,516.15,0,1,92679
563,1,0,1,1,59,1,1,Fiber optic,0,0,1,1,Two year,1,Credit card (automatic),99.5,5861.75,0,49,16,41.09,4583,0,Westminster,1,1,Fiber Optic,33.752590999999995,-117.99366100000002,1,99.5,1,3,None,88230,0,0,1,1,59,0,938.0,2424.3100000000004,0.0,5861.75,0,0,92683
564,1,0,0,0,7,1,0,DSL,0,0,1,0,Month-to-month,0,Bank transfer (automatic),64.3,445.95,0,19,58,31.84,4010,0,Rancho Santa Margarita,1,1,Fiber Optic,33.624654,-117.611733,0,64.3,0,0,Offer E,42193,1,2,0,0,7,1,259.0,222.88,0.0,445.95,1,0,92688
565,1,0,1,1,71,1,0,DSL,1,0,0,1,Two year,1,Credit card (automatic),70.85,4973.4,0,19,58,2.43,5328,0,Mission Viejo,1,1,DSL,33.611945,-117.66586699999999,1,70.85,0,3,None,46371,1,0,1,1,71,1,2885.0,172.53,0.0,4973.4,1,0,92691
566,1,0,1,1,15,1,0,Fiber optic,1,0,1,1,One year,0,Electronic check,101.9,1667.25,0,23,30,2.12,3707,0,Mission Viejo,0,1,Fiber Optic,33.60693,-117.644253,1,101.9,1,8,None,46227,1,1,1,1,15,2,0.0,31.8,0.0,1667.25,1,1,92692
567,1,0,1,0,71,1,1,DSL,1,1,1,0,Two year,0,Credit card (automatic),73.5,5357.75,0,34,5,34.39,5431,0,Ladera Ranch,0,1,DSL,33.569186,-117.640055,1,73.5,0,7,None,350,1,0,1,0,71,0,268.0,2441.69,0.0,5357.75,0,0,92694
568,0,0,0,0,35,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.25,3527.6,1,44,19,10.49,2744,1,Santa Ana,1,0,DSL,33.748478000000006,-117.85891799999999,0,104.26,0,0,Offer C,58157,0,1,0,1,35,2,670.0,367.15,0.0,3527.6,0,0,92701
569,0,0,0,0,11,0,No phone service,DSL,0,1,0,0,One year,1,Credit card (automatic),40.4,422.6,0,23,59,0.0,2133,0,Santa Ana,1,0,Cable,33.748635,-117.906125,0,40.4,0,0,None,70011,1,0,0,0,11,0,249.0,0.0,0.0,422.6,1,0,92703
570,0,0,1,1,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.25,1103.25,0,32,0,23.68,6134,0,Santa Ana,0,0,NA,33.719869,-117.907063,1,19.25,3,2,None,91188,0,0,1,0,60,0,0.0,1420.8,0.0,1103.25,0,0,92704
571,1,1,0,0,47,1,1,DSL,0,1,0,0,Two year,0,Bank transfer (automatic),59.6,2754,0,74,10,14.78,3155,0,Santa Ana,0,1,Fiber Optic,33.766003999999995,-117.786763,0,59.6,0,0,None,44117,1,0,0,0,47,0,0.0,694.66,0.0,2754.0,0,1,92705
572,0,0,0,0,11,1,0,DSL,0,0,0,1,One year,0,Credit card (automatic),64.9,697.25,0,55,23,5.0,3206,0,Santa Ana,1,0,Fiber Optic,33.765893,-117.881533,0,64.9,0,0,None,37879,1,0,0,1,11,0,0.0,55.0,0.0,697.25,0,1,92706
573,1,0,1,0,56,1,1,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),100.3,5614.45,1,50,8,26.15,5170,1,Santa Ana,0,1,Cable,33.714828999999995,-117.872941,1,104.31200000000001,0,2,None,62634,0,0,1,1,56,0,449.0,1464.4,0.0,5614.45,0,0,92707
574,0,1,1,0,28,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,110.85,3204.4,0,76,8,45.67,3906,0,Fountain Valley,1,0,DSL,33.712036,-117.95011299999999,1,110.85,0,6,Offer C,54548,1,0,1,0,28,0,0.0,1278.76,0.0,3204.4,0,1,92708
575,1,0,1,0,61,1,0,DSL,1,1,1,1,Two year,1,Mailed check,81.05,4747.65,0,26,51,20.34,4072,0,Tustin,0,1,Fiber Optic,33.735802,-117.818805,1,81.05,0,2,None,55062,1,0,1,1,61,1,0.0,1240.74,0.0,4747.65,1,1,92780
576,1,0,1,1,31,1,1,Fiber optic,1,0,1,0,One year,0,Bank transfer (automatic),98.05,3082.1,0,27,59,36.49,4524,0,Tustin,1,1,Fiber Optic,33.738543,-117.785046,1,98.05,3,3,Offer C,17494,0,0,1,0,31,2,0.0,1131.19,0.0,3082.1,1,1,92782
577,1,0,0,0,9,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.5,597.9,0,30,52,40.71,3198,0,Anaheim,0,1,Fiber Optic,33.844983,-117.952151,0,70.5,0,0,Offer E,60553,0,0,0,0,9,0,31.09,366.39,0.0,597.9,0,1,92801
578,1,1,1,0,35,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,94.55,3365.4,0,68,18,20.44,2631,0,Anaheim,0,1,Fiber Optic,33.807864,-117.923782,1,94.55,0,3,Offer C,45086,0,0,1,0,35,0,606.0,715.4000000000002,0.0,3365.4,0,0,92802
579,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.65,38.8,0,59,0,9.61,3007,0,Anaheim,0,1,NA,33.818000000000005,-117.974404,0,19.65,0,0,Offer E,81333,0,0,0,0,2,0,0.0,19.22,0.0,38.8,0,0,92804
580,0,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.0,233.55,1,48,0,19.48,3535,1,Anaheim,0,0,NA,33.830209,-117.906099,1,19.0,0,1,Offer D,68802,0,1,1,0,12,3,0.0,233.76,0.0,233.55,0,0,92805
581,0,0,0,0,1,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Mailed check,75.3,75.3,1,28,56,4.13,3244,1,Anaheim,0,0,Cable,33.837959999999995,-117.870494,0,78.312,0,0,None,34398,0,0,0,0,1,0,0.0,4.13,0.0,75.3,1,0,92806
582,0,1,0,0,4,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,89.2,346.2,1,74,26,48.35,5808,1,Anaheim,1,0,Cable,33.848733,-117.788357,0,92.76799999999999,0,0,None,36301,0,2,0,0,4,2,0.0,193.4,0.0,346.2,0,1,92807
583,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.0,19,0,62,0,28.28,2400,0,Anaheim,0,0,NA,33.850452000000004,-117.72666799999999,1,19.0,1,1,Offer E,19629,0,0,1,0,1,0,0.0,28.28,0.0,19.0,0,0,92808
584,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.0,61.7,0,40,0,15.37,5575,0,Brea,0,0,NA,33.930199,-117.862898,0,20.0,0,0,Offer E,34055,0,0,0,0,3,0,0.0,46.11,0.0,61.7,0,0,92821
585,0,1,0,0,1,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.7,85.7,1,68,23,45.81,4880,1,Brea,0,0,Cable,33.924143,-117.79387,0,89.12799999999999,0,0,None,1408,0,1,0,0,1,5,0.0,45.81,0.0,85.7,0,0,92823
586,1,0,0,0,52,1,0,DSL,1,1,1,0,Two year,1,Credit card (automatic),63.25,3342.45,0,56,10,46.24,6471,0,Fullerton,0,1,Fiber Optic,33.879983,-117.895482,0,63.25,0,0,None,34592,0,0,0,0,52,2,0.0,2404.48,0.0,3342.45,0,1,92831
587,1,0,1,1,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,85.1,0,28,0,5.2,2894,0,Fullerton,0,1,NA,33.868316,-117.929029,1,20.1,0,1,None,24502,0,0,1,0,5,0,0.0,26.0,0.0,85.1,1,0,92832
588,1,0,1,0,72,1,1,Fiber optic,1,1,0,1,Two year,1,Electronic check,99.15,7422.1,0,52,8,28.86,5152,0,Fullerton,1,1,DSL,33.877639,-117.96121200000002,1,99.15,0,1,None,46105,0,0,1,1,72,1,0.0,2077.92,0.0,7422.1,0,1,92833
589,1,0,1,1,71,1,1,DSL,1,1,1,1,Two year,0,Electronic check,90.4,6668.05,0,25,52,3.57,5633,0,Fullerton,1,1,DSL,33.902211,-117.914922,1,90.4,0,1,None,21157,1,0,1,1,71,0,0.0,253.47,0.0,6668.05,1,1,92835
590,1,0,1,0,72,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),111.9,8071.05,0,32,27,47.83,6437,0,Garden Grove,1,1,Fiber Optic,33.787165,-117.93188899999998,1,111.9,0,1,None,50641,1,0,1,1,72,3,0.0,3443.76,0.0,8071.05,0,1,92840
591,1,0,1,1,46,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,24.9,1174.8,0,56,0,18.45,2026,0,Garden Grove,0,1,NA,33.786738,-117.982564,1,24.9,0,1,None,31428,0,0,1,0,46,2,0.0,848.6999999999998,0.0,1174.8,0,0,92841
592,1,0,1,1,63,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),83.5,5435,0,19,69,13.45,4652,0,Garden Grove,1,1,Fiber Optic,33.764018,-117.93150700000001,1,83.5,0,1,None,43491,0,0,1,1,63,1,3750.0,847.3499999999998,0.0,5435.0,1,0,92843
593,1,0,0,0,30,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),84.3,2438.6,0,52,20,24.73,5393,0,Garden Grove,1,1,Cable,33.766476000000004,-117.96979499999999,0,84.3,0,0,Offer C,23481,0,0,0,0,30,0,0.0,741.9,0.0,2438.6,0,1,92844
594,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.6,45.6,0,36,9,37.44,2352,0,Garden Grove,0,1,Fiber Optic,33.782955,-118.02645600000001,0,45.6,0,0,None,15878,0,0,0,0,1,2,0.0,37.44,0.0,45.6,0,1,92845
595,0,0,0,0,12,1,1,DSL,1,0,0,0,Month-to-month,1,Mailed check,61.65,713.75,1,52,33,36.24,5670,1,Norco,1,0,Cable,33.925833000000004,-117.55963899999999,0,64.116,0,0,Offer D,22443,1,0,0,0,12,0,0.0,434.88,0.0,713.75,0,1,92860
596,1,0,0,0,16,0,No phone service,DSL,1,1,1,0,Two year,0,Mailed check,54.85,916.15,0,45,27,0.0,2136,0,Villa Park,1,1,Cable,33.817473,-117.81046200000002,0,54.85,0,0,None,5935,1,0,0,0,16,2,0.0,0.0,0.0,916.15,0,1,92861
597,1,0,0,0,4,1,1,DSL,0,0,0,1,Month-to-month,0,Mailed check,65.55,237.2,0,22,59,13.31,5707,0,Orange,0,1,Fiber Optic,33.828779,-117.848299,0,65.55,0,0,None,18058,1,0,0,1,4,0,140.0,53.24,0.0,237.2,1,0,92865
598,1,0,1,0,51,1,1,Fiber optic,0,1,0,1,One year,1,Credit card (automatic),90.35,4614.55,0,53,30,9.21,4965,0,Orange,0,1,DSL,33.784597,-117.84453500000001,1,90.35,0,0,None,15396,0,0,0,1,51,3,1384.0,469.71,0.0,4614.55,0,0,92866
599,1,0,1,0,65,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.4,1414.45,0,59,0,23.46,5368,0,Orange,0,1,NA,33.81859,-117.821288,1,20.4,0,1,None,40915,0,0,1,0,65,1,0.0,1524.9,0.0,1414.45,0,0,92867
600,1,0,0,0,16,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.55,1170.5,0,21,82,38.32,2893,0,Orange,0,1,Fiber Optic,33.787796,-117.875928,0,74.55,0,0,None,23172,1,0,0,0,16,1,960.0,613.12,0.0,1170.5,1,0,92868
601,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.95,47.7,0,47,0,31.45,3488,0,Orange,0,1,NA,33.792790999999994,-117.789749,0,19.95,0,0,None,37916,0,0,0,0,2,1,0.0,62.9,0.0,47.7,0,0,92869
602,0,0,1,1,66,1,1,Fiber optic,0,0,0,0,One year,1,Bank transfer (automatic),74.25,4859.25,0,34,17,37.84,4395,0,Placentia,0,0,Cable,33.881158,-117.85478300000001,1,74.25,1,1,None,48170,0,0,1,0,66,0,82.61,2497.44,0.0,4859.25,0,1,92870
603,1,0,0,0,46,1,1,Fiber optic,0,1,1,1,Two year,0,Electronic check,108.65,4903.2,0,51,22,37.5,4210,0,Corona,1,1,DSL,33.893823,-117.531446,0,108.65,0,0,None,44875,1,0,0,1,46,0,107.87,1725.0,0.0,4903.2,0,1,92879
604,0,0,0,0,32,1,1,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),109.55,3608,0,55,12,4.61,5076,0,Corona,1,0,DSL,33.918043,-117.61780900000001,0,109.55,0,0,None,16998,1,0,0,1,32,1,43.3,147.52,0.0,3608.0,0,1,92880
605,1,0,1,0,72,1,1,DSL,1,0,1,1,Two year,0,Credit card (automatic),86.65,6094.25,0,35,23,12.12,5483,0,Corona,1,1,Fiber Optic,33.833686,-117.51306299999999,1,86.65,0,1,None,21911,1,0,1,1,72,0,0.0,872.64,3.2,6094.25,0,1,92881
606,1,0,1,1,38,1,0,DSL,1,0,1,1,Two year,0,Credit card (automatic),81.0,3084.9,0,28,73,22.05,3067,0,Corona,1,1,Fiber Optic,33.819385,-117.60021299999998,1,81.0,0,1,None,60294,1,0,1,1,38,1,0.0,837.9,0.0,3084.9,1,1,92882
607,1,0,0,1,51,1,0,DSL,0,0,0,0,One year,0,Credit card (automatic),47.85,2356.75,0,48,20,36.59,4138,0,Corona,0,1,Fiber Optic,33.762351,-117.488725,0,47.85,0,0,None,13188,1,0,0,0,51,1,0.0,1866.09,18.39,2356.75,0,1,92883
608,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),114.55,8306.05,0,47,58,21.89,6158,0,Yorba Linda,1,1,Fiber Optic,33.897253000000006,-117.792202,1,114.55,3,1,None,39458,1,0,1,1,72,1,0.0,1576.08,21.6,8306.05,0,1,92886
609,0,1,1,0,65,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Bank transfer (automatic),105.25,6786.4,1,78,31,18.39,4196,1,Yorba Linda,1,0,Cable,33.884073,-117.732197,1,109.46,0,3,Offer B,20893,0,0,1,0,65,5,0.0,1195.35,0.0,6786.4,0,1,92887
610,1,0,1,1,9,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,29.95,248.95,1,32,10,0.0,2573,1,Ventura,0,1,Cable,34.360261,-119.30638300000001,1,31.148000000000003,0,1,Offer E,32899,0,0,1,0,9,2,0.0,0.0,0.0,248.95,0,1,93001
611,0,0,1,1,9,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,65.0,663.05,1,20,76,6.35,3983,1,Ventura,1,0,DSL,34.279221,-119.22143700000001,1,67.60000000000001,0,1,Offer E,46894,1,0,1,0,9,1,504.0,57.15,0.0,663.05,1,0,93003
612,1,0,0,1,66,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.55,1357.1,0,57,0,20.63,4101,0,Ventura,0,1,NA,34.278696999999994,-119.167798,0,20.55,2,0,None,27381,0,0,0,0,66,0,0.0,1361.58,17.14,1357.1,0,0,93004
613,0,1,0,0,44,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),109.8,4860.35,0,71,2,49.75,5720,0,Camarillo,1,0,Fiber Optic,34.227846,-119.079903,0,109.8,0,0,None,42853,0,0,0,0,44,0,0.0,2189.0,0.0,4860.35,0,1,93010
614,1,0,0,0,50,1,1,DSL,0,0,0,1,Two year,0,Bank transfer (automatic),69.5,3418.2,0,63,2,27.04,4145,0,Camarillo,1,1,Cable,34.205504,-118.99311100000001,0,69.5,0,0,None,24945,1,0,0,1,50,2,0.0,1352.0,5.73,3418.2,0,1,93012
615,0,0,0,0,15,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,48.85,631.4,0,64,19,13.58,3762,0,Carpinteria,0,0,DSL,34.441398,-119.51316299999999,0,48.85,0,0,None,17409,0,0,0,0,15,0,0.0,203.7,32.09,631.4,0,1,93013
616,1,0,0,0,8,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),25.25,186.3,0,55,16,0.0,2372,0,Fillmore,0,1,Fiber Optic,34.408161,-118.86511100000001,0,25.25,0,0,None,16013,0,0,0,0,8,0,30.0,0.0,0.0,186.3,0,0,93015
617,0,1,0,0,66,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),102.85,6976.75,0,69,5,11.63,5569,0,Moorpark,1,0,Fiber Optic,34.312945,-118.85816899999999,0,102.85,0,0,Offer A,32984,1,0,0,0,66,0,0.0,767.58,0.0,6976.75,0,1,93021
618,0,0,0,0,57,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Bank transfer (automatic),87.55,4884.85,0,30,41,28.27,4882,0,Oak View,0,0,Fiber Optic,34.404544,-119.302118,0,87.55,0,0,None,6503,1,2,0,0,57,3,0.0,1611.39,1.83,4884.85,0,1,93022
619,0,0,0,0,7,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),78.55,522.95,0,51,16,40.76,4025,0,Ojai,0,0,Fiber Optic,34.581308,-118.93194799999999,0,78.55,0,0,None,21633,0,0,0,0,7,1,0.0,285.32,47.19,522.95,0,1,93023
620,1,1,1,1,10,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Bank transfer (automatic),34.55,362.6,0,73,53,0.0,5248,0,Oxnard,0,1,DSL,34.223244,-119.18012,1,34.55,3,1,None,79736,0,0,1,0,10,2,0.0,0.0,0.0,362.6,0,1,93030
621,0,0,0,0,62,1,1,Fiber optic,1,1,0,0,One year,1,Electronic check,92.05,5755.8,0,27,47,23.88,5801,0,Oxnard,1,0,DSL,34.156628999999995,-119.117218,0,92.05,0,0,None,77791,0,0,0,0,62,0,2705.0,1480.56,14.21,5755.8,1,0,93033
622,1,0,1,1,40,1,0,Fiber optic,0,0,1,0,One year,1,Electronic check,85.05,3355.65,0,56,22,14.41,5904,0,Oxnard,1,1,Fiber Optic,34.184540000000005,-119.22466599999998,1,85.05,1,5,None,25322,0,0,1,0,40,0,0.0,576.4,38.15,3355.65,0,1,93035
623,0,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.7,406.95,0,49,0,15.87,4404,0,Piru,0,0,NA,34.432843,-118.730106,0,19.7,0,0,None,1459,0,0,0,0,20,2,0.0,317.4,0.0,406.95,0,0,93040
624,0,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.0,137.6,1,27,0,16.04,4479,1,Port Hueneme,0,0,NA,34.110124,-119.100972,0,20.0,0,0,Offer E,25634,0,0,0,0,7,3,0.0,112.28,0.0,137.6,1,0,93041
625,0,0,1,0,25,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.15,2395.7,0,22,52,29.81,3273,0,Santa Paula,0,0,Fiber Optic,34.402343,-119.094824,1,95.15,0,0,None,32511,1,0,0,1,25,1,0.0,745.25,0.0,2395.7,1,1,93060
626,1,0,1,0,23,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,84.25,1968.1,0,28,51,18.05,2781,0,Simi Valley,1,1,Fiber Optic,34.296813,-118.685703,1,84.25,0,1,None,49027,0,0,1,0,23,2,0.0,415.15,8.3,1968.1,1,1,93063
627,0,1,1,0,66,1,1,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),104.6,6819.45,0,74,15,25.51,5722,0,Simi Valley,1,0,DSL,34.269449,-118.76847099999999,1,104.6,0,7,Offer A,64802,0,0,1,0,66,1,1023.0,1683.66,0.0,6819.45,0,0,93065
628,0,1,0,0,72,1,1,Fiber optic,0,1,1,1,Two year,0,Electronic check,111.65,7943.45,0,72,14,44.81,5388,0,Somis,1,0,DSL,34.297628,-119.014627,0,111.65,0,0,Offer A,2966,1,1,0,0,72,1,0.0,3226.32,0.0,7943.45,0,1,93066
629,1,1,1,0,49,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Credit card (automatic),90.05,4547.25,1,75,15,22.92,5059,1,Summerland,0,1,Cable,34.420998,-119.60136999999999,1,93.652,0,3,Offer B,576,0,0,1,0,49,5,0.0,1123.0800000000004,0.0,4547.25,0,1,93067
630,1,1,1,1,43,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),110.75,4687.9,1,77,6,14.52,2728,1,Santa Barbara,1,1,DSL,34.419203,-119.710008,1,115.18,0,1,Offer B,31727,1,1,1,0,43,1,0.0,624.36,0.0,4687.9,0,1,93101
631,0,0,1,0,46,1,1,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),55.0,2473.95,0,48,15,13.05,5928,0,Santa Barbara,0,0,Fiber Optic,34.438581,-119.685368,1,55.0,0,9,None,20893,0,0,1,0,46,0,0.0,600.3000000000002,31.39,2473.95,0,1,93103
632,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.85,6562.9,0,41,9,26.96,6046,0,Santa Barbara,1,1,Fiber Optic,34.037341999999995,-119.80078999999999,1,89.85,0,5,None,25771,1,0,1,1,72,0,591.0,1941.12,12.55,6562.9,0,0,93105
633,1,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.35,176.3,0,40,0,17.4,4745,0,Santa Barbara,0,1,NA,34.457541,-119.631072,0,20.35,0,0,None,12741,0,0,0,0,10,0,0.0,174.0,0.0,176.3,0,0,93108
634,0,0,0,0,40,0,No phone service,DSL,1,0,1,1,One year,1,Bank transfer (automatic),54.55,2236.2,0,31,28,0.0,3533,0,Santa Barbara,0,0,DSL,34.406256,-119.72693600000001,0,54.55,0,0,Offer B,10986,1,0,0,1,40,2,626.0,0.0,11.48,2236.2,0,0,93109
635,0,0,1,1,65,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.5,6985.65,1,20,29,34.14,5720,1,Santa Barbara,1,0,Cable,34.437945,-119.77191,1,109.72,0,7,None,15757,0,3,1,1,65,4,2026.0,2219.1,0.0,6985.65,1,0,93110
636,1,0,0,0,31,1,0,Fiber optic,0,0,1,1,Two year,0,Bank transfer (automatic),99.45,3109.9,0,41,14,10.05,2021,0,Santa Barbara,1,1,Fiber Optic,34.460196999999994,-119.80260200000001,0,99.45,0,0,None,16477,1,0,0,1,31,0,435.0,311.55,43.38,3109.9,0,0,93111
637,0,0,1,0,68,1,1,DSL,1,1,0,0,Two year,0,Credit card (automatic),70.9,4911.35,0,48,9,27.41,4114,0,Goleta,1,0,DSL,34.489983,-120.091246,1,70.9,0,2,None,49975,1,0,1,0,68,0,0.0,1863.88,49.37,4911.35,0,1,93117
638,1,1,1,1,56,1,1,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),104.55,5794.65,1,80,13,48.8,6268,1,Alpaugh,1,1,DSL,35.869626000000004,-119.49877099999999,1,108.73200000000001,0,0,Offer B,1054,0,0,0,0,56,0,753.0,2732.8,0.0,5794.65,0,0,93201
639,1,0,1,0,10,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.25,855.3,1,26,90,2.02,3573,1,Armona,0,1,DSL,36.315979,-119.710852,1,88.66,0,1,Offer D,2872,0,0,1,1,10,0,770.0,20.2,0.0,855.3,1,0,93202
640,1,0,1,1,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.4,1620.2,0,50,0,19.09,5668,0,Arvin,0,1,NA,35.116307,-118.817644,1,25.4,2,10,None,16206,0,0,1,0,68,1,0.0,1298.12,9.34,1620.2,0,0,93203
641,0,0,1,1,43,1,0,DSL,0,0,1,0,Month-to-month,0,Electronic check,56.15,2499.3,1,57,22,37.25,2152,1,Avenal,0,0,Cable,35.916942999999996,-120.129921,1,58.396,0,3,None,14697,0,1,1,0,43,6,550.0,1601.75,0.0,2499.3,0,0,93204
642,1,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.55,89.55,1,38,30,42.46,4996,1,Bodfish,0,1,Fiber Optic,35.523990999999995,-118.40043200000001,0,93.132,0,0,Offer E,1954,0,3,0,1,1,2,0.0,42.46,0.0,89.55,0,1,93205
643,0,1,0,0,49,1,0,Fiber optic,0,1,0,1,One year,1,Bank transfer (automatic),89.85,4287.2,0,70,21,47.72,5982,0,Buttonwillow,1,0,Cable,35.451402,-119.488413,0,89.85,0,0,None,2078,0,0,0,0,49,0,0.0,2338.28,0.0,4287.2,0,1,93206
644,0,0,1,1,15,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,25.25,394.85,0,21,0,29.55,4667,0,California Hot Springs,0,0,NA,35.865795,-118.69758999999999,1,25.25,1,1,None,226,0,0,1,0,15,1,0.0,443.25,0.0,394.85,1,0,93207
645,1,1,1,0,20,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.55,1899.65,1,75,11,5.31,5604,1,Camp Nelson,0,1,Cable,36.057458000000004,-118.591951,1,98.33200000000001,0,7,None,191,0,3,1,1,20,2,209.0,106.2,0.0,1899.65,0,0,93208
646,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.7,45.7,1,57,14,5.55,2295,1,Coalinga,0,1,Fiber Optic,36.186867,-120.38779299999999,0,47.52800000000001,0,0,Offer E,18036,0,1,0,0,1,2,0.0,5.55,0.0,45.7,0,0,93210
647,1,0,1,1,50,1,1,DSL,0,0,1,0,One year,1,Electronic check,69.65,3442.15,0,25,58,14.32,4706,0,Corcoran,1,1,DSL,36.04533,-119.532424,1,69.65,0,6,Offer B,23506,1,0,1,0,50,1,1996.0,716.0,0.0,3442.15,1,0,93212
648,0,1,0,0,2,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,89.5,161.5,1,69,21,47.47,2065,1,Delano,0,0,DSL,35.772244,-119.20968899999998,0,93.08,0,0,None,37280,0,0,0,1,2,5,34.0,94.94,0.0,161.5,0,0,93215
649,1,1,0,0,24,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),70.0,1732.6,0,74,13,31.73,5242,0,Ducor,0,1,DSL,35.846067,-119.00407299999999,0,70.0,0,0,Offer C,823,0,0,0,0,24,0,0.0,761.52,0.0,1732.6,0,1,93218
650,0,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.55,222.3,1,30,33,26.26,2876,1,Earlimart,0,0,Fiber Optic,35.858053999999996,-119.305858,0,72.332,0,0,None,9318,0,2,0,0,3,2,7.34,78.78,0.0,222.3,0,1,93219
651,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.6,74.6,1,23,52,22.16,3860,1,Exeter,1,0,Fiber Optic,36.301689,-119.01823300000001,0,77.584,0,0,Offer E,13333,0,0,0,0,1,4,0.0,22.16,0.0,74.6,1,0,93221
652,1,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.1,655.3,0,37,0,11.75,4517,0,Frazier Park,0,1,NA,34.907911,-119.23428100000001,1,20.1,3,7,None,1526,0,0,1,0,35,2,0.0,411.25,38.61,655.3,0,0,93222
653,0,0,0,0,17,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,24.8,475.25,0,64,0,9.84,5208,0,Farmersville,0,0,NA,36.29878,-119.20102800000001,0,24.8,0,0,Offer D,8644,0,0,0,0,17,0,0.0,167.28,37.06,475.25,0,0,93223
654,0,1,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.65,164.3,1,74,0,27.95,5432,1,Fellows,0,0,NA,35.215731,-119.57013,0,19.65,0,0,None,626,0,0,0,0,8,6,0.0,223.6,0.0,164.3,0,0,93224
655,1,0,0,0,10,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),95.1,865.1,0,32,11,45.69,5787,0,Frazier Park,0,1,Fiber Optic,34.827662,-118.999073,0,95.1,0,0,Offer D,4498,1,0,0,1,10,0,95.0,456.9,43.25,865.1,0,0,93225
656,1,0,1,1,68,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),88.85,6132.7,0,39,14,41.61,5228,0,Glennville,1,1,Fiber Optic,35.735694,-118.738483,1,88.85,0,2,None,296,1,0,1,1,68,0,859.0,2829.48,0.0,6132.7,0,0,93226
657,1,0,1,0,45,1,0,DSL,1,1,1,1,One year,0,Bank transfer (automatic),78.8,3597.5,0,38,19,9.91,4192,0,Hanford,1,1,Cable,36.292229999999996,-119.622676,1,78.8,0,6,Offer B,53204,0,0,1,1,45,0,684.0,445.95,23.28,3597.5,0,0,93230
658,1,0,1,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.85,35.9,1,40,0,15.14,2362,1,Huron,0,1,NA,36.217864,-120.08011699999999,1,19.85,0,2,Offer E,6918,0,1,1,0,2,4,0.0,30.28,0.0,35.9,0,0,93234
659,1,0,1,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.35,697.65,0,56,0,2.15,3078,0,Ivanhoe,0,1,NA,36.385818,-119.22424299999999,1,20.35,0,3,None,4517,0,0,1,0,37,0,0.0,79.55,45.07,697.65,0,0,93235
660,0,0,0,0,4,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,24.25,96.05,1,48,18,0.0,2038,1,Kernville,0,0,Fiber Optic,35.852892,-118.397782,0,25.22,0,0,Offer E,1873,0,0,0,0,4,1,17.0,0.0,0.0,96.05,0,0,93238
661,0,0,0,0,10,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.25,428.7,0,46,29,3.55,5369,0,Kettleman City,0,0,Fiber Optic,35.996922999999995,-120.000951,0,45.25,0,0,Offer D,1809,0,0,0,0,10,1,12.43,35.5,44.9,428.7,0,1,93239
662,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,20.05,0,23,0,18.15,2798,0,Lake Isabella,0,1,NA,35.607875,-118.46631799999999,0,20.05,0,0,None,5564,0,0,0,0,1,0,0.0,18.15,0.0,20.05,1,0,93240
663,1,0,1,1,65,1,1,DSL,1,1,0,1,Two year,1,Mailed check,69.55,4459.15,0,40,30,17.43,5420,0,Lamont,0,1,Fiber Optic,35.245034999999994,-118.905553,1,69.55,0,10,Offer B,15364,0,0,1,1,65,0,133.77,1132.95,23.61,4459.15,0,1,93241
664,0,0,1,1,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.5,1167.6,0,33,0,42.14,5864,0,Laton,0,0,NA,36.444232,-119.71828500000001,1,19.5,3,5,Offer B,2900,0,0,1,0,57,0,0.0,2401.98,19.89,1167.6,0,0,93242
665,0,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.75,238.1,0,48,4,12.5,3319,0,Lebec,1,0,Fiber Optic,34.845861,-118.88516299999999,0,74.75,0,0,None,1247,0,0,0,0,3,0,0.95,37.5,38.84,238.1,0,1,93243
666,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.65,145.15,1,52,30,7.64,2323,1,Lemon Cove,0,0,Cable,36.462671,-118.99729099999999,0,72.436,0,0,Offer E,293,0,1,0,0,2,3,44.0,15.28,0.0,145.15,0,0,93244
667,1,0,0,0,49,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),30.2,1453.1,0,22,58,0.0,5214,0,Lemoore,1,1,Cable,36.303666,-119.825657,0,30.2,0,0,Offer B,30419,0,0,0,0,49,2,0.0,0.0,0.0,1453.1,1,1,93245
668,0,0,0,0,4,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.65,191.05,1,47,30,45.4,2864,1,Lindsay,0,0,Cable,36.205465000000004,-119.085807,0,47.476000000000006,0,0,None,15508,0,1,0,0,4,4,57.0,181.6,0.0,191.05,0,0,93247
669,0,0,1,0,70,0,No phone service,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),57.8,4039.3,0,22,85,0.0,5640,0,Lost Hills,1,0,Fiber Optic,35.637715,-119.893068,1,57.8,0,9,None,2502,1,0,1,1,70,2,0.0,0.0,1.01,4039.3,1,1,93249
670,0,0,1,1,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.85,1039.45,0,60,0,11.35,4836,0,Mc Farland,0,0,NA,35.666886,-119.18671699999999,1,19.85,0,6,Offer B,10781,0,0,1,0,53,0,0.0,601.55,14.67,1039.45,0,0,93250
671,1,0,1,1,53,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.55,1336.1,0,37,0,33.31,5794,0,Mc Kittrick,0,1,NA,35.38381,-119.73088500000001,1,25.55,3,3,Offer B,302,0,0,1,0,53,3,0.0,1765.43,37.37,1336.1,0,0,93251
672,0,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,75.05,75.05,1,23,64,32.86,4838,1,Temecula,0,0,DSL,33.507255,-117.029473,0,78.05199999999999,0,0,Offer E,46171,0,0,0,0,1,8,0.0,32.86,0.0,75.05,1,0,92592
673,1,0,0,0,22,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),24.85,493.4,0,49,0,22.97,3534,0,New Cuyama,0,1,NA,34.956577,-119.750142,0,24.85,0,0,Offer D,798,0,0,0,0,22,1,0.0,505.34,21.32,493.4,0,0,93254
674,1,1,0,0,52,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,49.15,2550.9,1,76,20,0.0,5597,1,Temecula,0,1,Cable,33.507255,-117.029473,0,51.11600000000001,0,0,None,46171,0,1,0,1,52,1,0.0,0.0,0.0,2550.9,0,1,92592
675,1,1,0,0,65,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,110.35,7246.15,0,80,27,44.23,4295,0,Pixley,1,1,DSL,35.957019,-119.330928,0,110.35,0,0,None,4198,1,0,0,0,65,1,0.0,2874.95,0.0,7246.15,0,1,93256
676,0,0,0,0,48,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),24.55,1203.95,0,63,0,23.76,5517,0,Porterville,0,0,NA,36.008958,-118.891593,0,24.55,0,0,Offer B,65566,0,0,0,0,48,0,0.0,1140.48,36.04,1203.95,0,0,93257
677,0,0,0,0,2,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,34.7,62.25,1,19,84,0.0,3146,1,Posey,0,0,Cable,35.861928000000006,-118.636698,0,36.088,0,0,Offer E,266,0,0,0,1,2,3,52.0,0.0,0.0,62.25,1,0,93260
678,1,0,0,0,3,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Mailed check,107.95,313.6,0,57,22,47.5,3449,0,Richgrove,1,1,Fiber Optic,35.809921,-119.12743700000001,0,107.95,0,0,None,2956,0,0,0,1,3,0,69.0,142.5,0.0,313.6,0,0,93261
679,1,0,1,0,45,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),81.4,3775.85,0,64,19,1.59,5602,0,Sequoia National Park,0,1,Fiber Optic,36.527243,-118.59493799999998,1,81.4,0,4,Offer B,56,0,0,1,0,45,1,0.0,71.55,0.0,3775.85,0,1,93262
680,1,0,1,1,1,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,80.0,80,1,48,3,35.71,2046,1,Shafter,0,1,Fiber Optic,35.490705,-119.286833,1,83.2,0,1,Offer E,15177,0,3,1,1,1,3,0.0,35.71,0.0,80.0,0,0,93263
681,0,0,1,1,61,1,0,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),73.8,4616.05,0,57,24,1.27,6301,0,Springville,1,0,DSL,36.245926000000004,-118.69313799999999,1,73.8,0,9,Offer B,3546,1,0,1,1,61,0,1108.0,77.47,49.51,4616.05,0,0,93265
682,1,0,0,0,3,1,0,DSL,1,0,1,0,Month-to-month,1,Credit card (automatic),64.4,195.65,0,37,7,38.05,5645,0,Stratford,0,1,Fiber Optic,36.175255,-119.813805,0,64.4,0,0,None,1729,1,0,0,0,3,0,1.37,114.15,0.0,195.65,0,1,93266
683,0,1,0,0,40,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),103.75,4188.4,0,74,24,28.54,3568,0,Strathmore,1,0,Cable,36.141319,-119.129075,0,103.75,0,0,None,5689,1,0,0,0,40,0,100.52,1141.6,0.0,4188.4,0,1,93267
684,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,71.1,71.1,0,47,10,37.51,3029,0,Taft,0,0,DSL,35.184837,-119.402525,0,71.1,0,0,None,14937,0,0,0,0,1,0,0.0,37.51,0.0,71.1,0,0,93268
685,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.9,49.9,0,33,4,14.93,4667,0,Terra Bella,0,0,Fiber Optic,35.939068,-119.04366599999999,0,49.9,0,0,None,5868,1,0,0,0,1,0,0.0,14.93,0.0,49.9,0,0,93270
686,1,0,0,0,51,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),24.6,1266.4,0,58,0,34.36,4886,0,Three Rivers,0,1,NA,36.413433000000005,-118.854708,0,24.6,0,0,Offer B,2318,0,0,0,0,51,0,0.0,1752.36,47.91,1266.4,0,0,93271
687,1,1,0,0,2,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.25,91.1,1,69,30,43.99,3475,1,San Diego,0,1,Fiber Optic,32.961064,-117.13491699999999,0,51.22,0,0,None,47224,0,0,0,0,2,5,27.0,87.98,0.0,91.1,0,0,92129
688,1,0,0,0,52,0,No phone service,DSL,0,1,0,0,One year,0,Mailed check,30.1,1623.4,0,42,14,0.0,6290,0,Tulare,0,1,DSL,36.185471,-119.375243,0,30.1,0,0,Offer B,56101,0,0,0,0,52,0,0.0,0.0,11.72,1623.4,0,1,93274
689,1,0,0,0,51,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Bank transfer (automatic),83.4,4149.45,0,55,12,45.92,4191,0,Tupman,0,1,DSL,35.316263,-119.40255900000001,0,83.4,0,0,Offer B,236,0,0,0,1,51,3,498.0,2341.92,29.76,4149.45,0,0,93276
690,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.45,20.45,0,53,0,11.61,5384,0,Visalia,0,1,NA,36.303793,-119.375646,0,20.45,0,0,None,44741,0,0,0,0,1,1,0.0,11.61,0.0,20.45,0,0,93277
691,1,0,1,1,31,1,1,DSL,1,1,0,1,One year,1,Bank transfer (automatic),75.25,2344.5,0,55,22,29.06,4258,0,Wasco,0,1,Cable,35.652242,-119.4464,1,75.25,0,7,None,22760,1,0,1,1,31,1,516.0,900.86,1.99,2344.5,0,0,93280
692,1,0,0,1,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.55,1013.05,0,62,0,42.25,3313,0,Weldon,0,1,NA,35.556470000000004,-118.244914,0,20.55,0,0,Offer B,1935,0,0,0,0,47,2,0.0,1985.75,0.0,1013.05,0,0,93283
693,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.1,270.7,1,63,11,26.52,4965,1,San Diego,0,0,DSL,32.961064,-117.13491699999999,0,78.104,0,0,Offer E,47224,0,1,0,0,3,6,30.0,79.56,0.0,270.7,0,0,92129
694,0,1,0,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.05,417,0,65,0,34.39,4327,0,Woodlake,0,0,NA,36.464634999999994,-119.094348,0,20.05,0,0,None,8870,0,0,0,0,22,0,0.0,756.58,0.0,417.0,0,0,93286
695,0,0,1,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.65,20.65,0,64,0,35.24,4517,0,Woody,0,0,NA,35.710244,-118.881679,1,20.65,0,8,None,88,0,0,1,0,1,0,0.0,35.24,0.0,20.65,0,0,93287
696,1,0,1,0,72,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),85.15,6316.2,0,19,52,32.36,6322,0,Visalia,1,1,DSL,36.391777000000005,-119.37284199999999,1,85.15,0,5,None,36718,1,0,1,1,72,0,3284.0,2329.92,0.0,6316.2,1,0,93291
697,1,0,1,1,3,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.15,168.15,1,23,56,13.54,3273,1,San Diego,1,1,Cable,32.961064,-117.13491699999999,1,52.156000000000006,0,1,None,47224,0,0,1,0,3,2,0.0,40.62,0.0,168.15,1,1,92129
698,1,1,1,1,47,1,0,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),84.95,4018.05,0,72,22,42.29,3384,0,Bakersfield,0,1,Fiber Optic,35.383937,-119.02042800000001,1,84.95,1,1,None,12963,0,1,1,0,47,3,884.0,1987.63,0.0,4018.05,0,0,93301
699,1,0,1,1,72,1,1,DSL,1,0,0,0,Two year,1,Credit card (automatic),66.5,4811.6,0,23,41,6.09,4397,0,Bakersfield,1,1,Cable,35.339796,-119.023552,1,66.5,0,8,None,44588,1,1,1,0,72,2,197.28,438.48,45.61,4811.6,1,1,93304
700,1,0,1,1,66,1,1,DSL,0,0,1,0,Two year,1,Bank transfer (automatic),63.3,4189.7,0,34,19,32.04,4186,0,Bakersfield,1,1,DSL,35.391733,-118.984109,1,63.3,0,5,None,35643,0,0,1,0,66,0,796.0,2114.64,40.62,4189.7,0,0,93305
701,1,0,0,0,35,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,83.15,2848.45,0,52,6,41.21,2332,0,Bakersfield,0,1,Fiber Optic,35.449881,-118.84144199999999,0,83.15,0,0,None,53481,0,0,0,0,35,0,171.0,1442.35,18.84,2848.45,0,0,93306
702,1,0,0,0,29,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.9,2516.2,0,56,21,9.49,4388,0,Bakersfield,0,1,Cable,35.280113,-118.962329,0,84.9,0,0,None,59195,0,0,0,1,29,0,0.0,275.21,47.04,2516.2,0,1,93307
703,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.55,33.6,0,30,0,16.7,5629,0,Bakersfield,0,0,NA,35.559616999999996,-118.92518500000001,0,20.55,0,0,None,44915,0,1,0,0,2,2,0.0,33.4,0.0,33.6,0,0,93308
704,1,0,0,0,4,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,49.25,208.45,0,34,5,38.01,3272,0,Bakersfield,0,1,Fiber Optic,35.342890999999995,-119.064803,0,49.25,0,0,None,58632,0,0,0,0,4,2,10.0,152.04,0.0,208.45,0,0,93309
705,0,0,0,0,25,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Bank transfer (automatic),79.85,2015.35,1,54,13,26.81,4535,1,San Diego,0,0,Fiber Optic,32.961064,-117.13491699999999,0,83.044,0,0,Offer C,47224,0,0,0,0,25,2,262.0,670.25,0.0,2015.35,0,0,92129
706,0,0,0,0,65,1,0,DSL,1,1,0,0,Two year,1,Mailed check,59.6,3739.8,0,19,76,43.29,4372,0,Bakersfield,0,0,DSL,35.392599,-119.245341,0,59.6,0,0,Offer B,40836,1,0,0,0,65,0,0.0,2813.85,0.0,3739.8,1,1,93312
707,1,1,0,0,27,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),104.65,2964,0,76,19,34.39,3104,0,Bakersfield,0,1,DSL,35.140938,-119.051348,0,104.65,0,0,Offer C,25126,1,0,0,0,27,3,0.0,928.53,0.0,2964.0,0,1,93313
708,1,0,1,0,29,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.3,2263.4,0,26,59,3.35,4910,0,San Luis Obispo,1,1,DSL,35.233745,-120.626442,1,75.3,0,10,None,27047,0,0,1,0,29,2,1335.0,97.15,0.0,2263.4,1,0,93401
709,1,0,1,1,29,1,1,DSL,0,1,1,1,Month-to-month,0,Credit card (automatic),80.1,2211.8,0,60,27,6.73,4558,0,Los Osos,1,1,Fiber Optic,35.279984000000006,-120.824288,1,80.1,2,6,None,14859,0,0,1,1,29,0,0.0,195.17,0.0,2211.8,0,1,93402
710,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.55,19.55,1,27,0,38.44,3556,1,San Diego,0,1,NA,32.961064,-117.13491699999999,0,19.55,0,0,None,47224,0,0,0,0,1,3,0.0,38.44,0.0,19.55,1,0,92129
711,0,0,1,0,20,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,81.0,1683.7,0,45,21,11.39,4741,0,Arroyo Grande,1,0,DSL,35.176235999999996,-120.48324299999999,1,81.0,0,6,Offer D,24499,1,0,1,0,20,2,354.0,227.8,0.0,1683.7,0,0,93420
712,0,0,0,0,58,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.7,1519,0,23,0,47.9,5138,0,Atascadero,0,0,NA,35.453912,-120.69461000000001,0,24.7,0,0,Offer B,29539,0,0,0,0,58,1,0.0,2778.2,0.0,1519.0,1,0,93422
713,0,0,0,1,14,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,86.0,1164.05,0,53,22,47.72,5494,0,Avila Beach,0,0,Fiber Optic,35.186644,-120.728305,0,86.0,1,0,Offer D,812,1,0,0,0,14,1,0.0,668.0799999999998,0.0,1164.05,0,1,93424
714,1,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.4,1710.9,0,61,0,34.29,5512,0,Bradley,0,1,NA,35.842889,-121.00486200000002,1,25.4,0,2,Offer A,1363,0,0,1,0,72,0,0.0,2468.88,0.0,1710.9,0,0,93426
715,1,0,0,0,46,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Credit card (automatic),89.15,4245.55,0,21,73,37.75,5593,0,Buellton,0,1,Fiber Optic,34.631362,-120.23821799999999,0,89.15,0,0,Offer B,4644,0,0,0,0,46,2,3099.0,1736.5,0.0,4245.55,1,0,93427
716,0,0,1,0,71,0,No phone service,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),58.25,4145.9,0,40,29,0.0,5224,0,Cambria,1,0,DSL,35.591387,-121.032256,1,58.25,0,2,Offer A,6526,1,0,1,1,71,0,1202.0,0.0,0.0,4145.9,0,0,93428
717,1,0,0,0,32,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),85.65,2664.3,0,51,28,37.04,2383,0,Casmalia,0,1,Cable,34.866032000000004,-120.536546,0,85.65,0,0,None,210,0,0,0,1,32,1,0.0,1185.28,0.0,2664.3,0,1,93429
718,0,0,0,0,26,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),50.35,1277.5,0,47,7,0.0,2510,0,Cayucos,1,0,DSL,35.511833,-120.91871299999998,0,50.35,0,0,None,3220,0,0,0,1,26,0,89.0,0.0,0.0,1277.5,0,0,93430
719,1,1,1,0,68,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),80.35,5589.3,0,75,15,34.31,5581,0,Creston,1,1,Fiber Optic,35.480896,-120.469476,1,80.35,0,7,Offer A,1203,0,0,1,0,68,0,838.0,2333.08,0.0,5589.3,0,0,93432
720,1,0,1,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.2,34.75,0,22,0,38.41,3866,0,Grover Beach,0,1,NA,35.120833000000005,-120.61843,1,20.2,0,6,None,13106,0,1,1,0,2,3,0.0,76.82,0.0,34.75,1,0,93433
721,1,0,1,1,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.55,1305.95,0,24,0,46.76,4446,0,Guadalupe,0,1,NA,34.936,-120.594655,1,20.55,0,0,Offer B,5726,0,0,0,0,61,0,0.0,2852.36,0.0,1305.95,1,0,93434
722,0,0,1,1,4,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.95,381.3,1,48,33,4.14,5640,1,San Diego,0,0,Fiber Optic,32.961064,-117.13491699999999,1,89.38799999999999,0,1,None,47224,0,0,1,1,4,2,12.58,16.56,0.0,381.3,0,1,92129
723,1,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.35,141.5,1,26,65,36.48,2450,1,San Diego,0,1,Cable,32.961064,-117.13491699999999,0,47.163999999999994,0,0,None,47224,0,0,0,0,3,5,92.0,109.44,0.0,141.5,1,0,92129
724,1,1,1,0,33,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.5,3105.55,1,72,9,27.78,4333,1,San Diego,0,1,Fiber Optic,32.961064,-117.13491699999999,1,98.28,0,1,None,47224,0,2,1,0,33,2,279.0,916.74,0.0,3105.55,0,0,92129
725,1,1,1,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,21.25,204.55,0,70,0,1.66,2302,0,Los Olivos,0,1,NA,34.70434,-120.02609,1,21.25,0,1,None,1317,0,0,1,0,9,0,0.0,14.94,0.0,204.55,0,0,93441
726,0,0,0,0,22,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,26.25,605.9,0,47,0,5.28,5676,0,Morro Bay,0,0,NA,35.369553,-120.76386399999998,0,26.25,0,0,Offer D,10909,0,0,0,0,22,1,0.0,116.16,0.0,605.9,0,0,93442
727,0,0,1,1,5,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.85,356.1,0,20,73,47.91,5109,0,Nipomo,0,0,Fiber Optic,35.050345,-120.489599,1,80.85,2,8,None,15405,0,0,1,0,5,0,26.0,239.55,0.0,356.1,1,1,93444
728,0,1,0,0,30,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Credit card (automatic),91.7,2758.15,1,69,21,45.88,2482,1,San Diego,1,0,Cable,32.961064,-117.13491699999999,0,95.368,0,0,None,47224,0,1,0,0,30,4,579.0,1376.4,0.0,2758.15,0,0,92129
729,1,0,0,0,65,1,1,DSL,0,1,0,1,Two year,1,Credit card (automatic),74.2,4805.65,0,41,18,22.23,4774,0,Paso Robles,1,1,Fiber Optic,35.634221999999994,-120.72834099999999,0,74.2,0,0,Offer B,35586,1,0,0,1,65,0,0.0,1444.95,0.0,4805.65,0,1,93446
730,0,0,0,0,45,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,87.25,3941.7,1,29,56,4.48,5269,1,San Diego,1,0,Cable,32.961064,-117.13491699999999,0,90.74,0,0,None,47224,1,0,0,0,45,2,2207.0,201.6,0.0,3941.7,1,0,92129
731,1,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,92.75,0,46,0,31.78,2303,0,San Ardo,0,1,NA,35.996008,-120.85305,0,20.35,0,0,None,670,0,0,0,0,5,0,0.0,158.9,0.0,92.75,0,0,93450
732,1,0,1,1,25,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,75.5,1901.05,0,51,58,4.46,5985,0,San Miguel,0,1,DSL,35.886767,-120.60866100000001,1,75.5,3,4,None,2666,0,0,1,0,25,1,110.26,111.5,0.0,1901.05,0,1,93451
733,0,0,1,1,72,1,1,Fiber optic,1,0,0,0,Two year,0,Bank transfer (automatic),79.05,5730.7,0,27,53,7.29,4689,0,San Simeon,0,0,Fiber Optic,35.746484,-121.223355,1,79.05,0,5,Offer A,471,0,0,1,0,72,1,0.0,524.88,0.0,5730.7,1,1,93452
734,0,0,1,0,27,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Bank transfer (automatic),90.15,2423.4,0,25,59,18.74,5750,0,Santa Margarita,1,0,Fiber Optic,35.303926000000004,-120.25656699999999,1,90.15,0,1,None,2687,0,0,1,1,27,2,0.0,505.98,0.0,2423.4,1,1,93453
735,1,0,1,1,32,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Credit card (automatic),50.6,1653.45,0,48,19,0.0,3087,0,Santa Maria,1,1,DSL,34.943523,-120.256729,1,50.6,2,10,None,30540,0,0,1,1,32,0,0.0,0.0,0.0,1653.45,0,1,93454
736,0,0,0,0,30,1,1,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),110.45,3327.05,0,19,27,13.16,4983,0,Santa Maria,1,0,Cable,34.818227,-120.418784,0,110.45,0,0,None,37364,1,0,0,1,30,0,0.0,394.8,0.0,3327.05,1,1,93455
737,1,0,1,0,70,1,0,Fiber optic,1,1,0,1,Two year,0,Credit card (automatic),101.0,7085.5,0,26,59,41.05,5025,0,Santa Maria,1,1,Fiber Optic,34.959340000000005,-120.490081,1,101.0,0,9,Offer A,43684,1,0,1,1,70,3,4180.0,2873.5,0.0,7085.5,1,0,93458
738,1,1,0,0,42,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),79.35,3344.1,0,66,19,13.51,2399,0,Santa Ynez,0,1,Fiber Optic,34.630356,-120.032564,0,79.35,0,0,None,5710,0,0,0,0,42,0,635.0,567.42,0.0,3344.1,0,0,93460
739,0,1,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),89.85,6697.35,0,68,17,48.51,5881,0,Shandon,1,0,Fiber Optic,35.634488,-120.29353400000001,1,89.85,0,0,Offer A,1255,1,0,0,0,72,0,0.0,3492.72,0.0,6697.35,0,1,93461
740,0,0,0,0,47,1,1,DSL,1,0,0,0,Two year,1,Mailed check,65.0,2879.9,0,38,13,35.75,3286,0,Solvang,1,0,DSL,34.624399,-120.137875,0,65.0,0,0,Offer B,7958,1,0,0,0,47,0,0.0,1680.25,0.0,2879.9,0,1,93463
741,0,0,0,0,2,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,80.45,137.1,0,35,25,35.41,5602,0,Templeton,1,0,Fiber Optic,35.536115,-120.739231,0,80.45,0,0,None,7918,0,0,0,0,2,0,34.0,70.82,0.0,137.1,0,0,93465
742,1,0,0,0,10,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Electronic check,98.55,1008.55,1,51,14,27.57,3658,1,San Diego,0,1,DSL,32.961064,-117.13491699999999,0,102.492,0,0,Offer D,47224,0,0,0,1,10,4,0.0,275.7,0.0,1008.55,0,1,92129
743,0,0,1,1,61,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.1,1551.6,0,23,0,13.35,5970,0,California City,0,0,NA,35.151491,-117.92759699999999,1,24.1,0,9,Offer B,8316,0,0,1,0,61,1,0.0,814.35,0.0,1551.6,1,0,93505
744,0,0,0,0,5,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),44.05,202.15,0,46,29,10.99,5846,0,Acton,0,0,Fiber Optic,34.501452,-118.207862,0,44.05,0,0,None,7831,0,0,0,0,5,0,59.0,54.95,0.0,202.15,0,0,93510
745,0,1,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),110.8,7882.25,0,69,2,15.85,5933,0,Benton,1,0,DSL,37.653946999999995,-118.231443,1,110.8,0,8,Offer A,340,1,0,1,0,72,0,158.0,1141.2,0.0,7882.25,0,0,93512
746,1,1,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.95,8196.4,0,75,2,21.38,6268,0,Big Pine,1,1,Cable,37.245505,-118.06294299999999,1,114.95,0,3,Offer A,1826,1,1,1,0,72,2,0.0,1539.36,0.0,8196.4,0,1,93513
747,0,1,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,75.05,202.9,0,74,13,41.44,3545,0,Bishop,1,0,Fiber Optic,37.045840000000005,-118.397236,0,75.05,0,0,Offer E,13309,0,0,0,0,3,0,0.0,124.32,5.49,202.9,0,1,93514
748,1,0,1,0,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.25,855.1,0,43,0,15.95,2282,0,Boron,0,1,NA,34.957029999999996,-117.73045,1,19.25,0,5,Offer B,2241,0,0,1,0,48,3,0.0,765.5999999999998,0.0,855.1,0,0,93516
749,0,0,0,0,63,1,0,Fiber optic,0,0,1,0,One year,1,Credit card (automatic),90.05,5817,0,41,8,40.34,4039,0,Bridgeport,1,0,Cable,38.184583,-119.28655800000001,0,90.05,0,0,Offer B,826,1,1,0,0,63,2,465.0,2541.42,0.0,5817.0,0,0,93517
750,0,0,0,0,27,1,0,DSL,1,1,0,0,Month-to-month,1,Mailed check,56.7,1652.95,0,35,9,25.21,4472,0,Caliente,0,0,Fiber Optic,35.358953,-118.527064,0,56.7,0,0,None,1022,0,0,0,0,27,0,0.0,680.6700000000002,0.0,1652.95,0,1,93518
751,1,0,1,1,70,1,0,DSL,1,1,1,1,Two year,1,Credit card (automatic),80.15,5600.15,0,28,46,24.08,5715,0,Darwin,1,1,Fiber Optic,36.319181,-117.593053,1,80.15,0,10,Offer A,64,0,2,1,1,70,1,257.61,1685.6,0.0,5600.15,1,1,93522
752,1,0,1,1,7,1,0,DSL,1,0,0,1,Month-to-month,1,Credit card (automatic),71.35,515.75,0,47,25,49.98,3459,0,Edwards,1,1,DSL,34.966777,-117.961179,1,71.35,2,3,None,7685,1,0,1,1,7,2,129.0,349.86,0.0,515.75,0,0,93523
753,1,0,0,1,0,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.25, ,0,24,0,13.16,5504,0,Independence,0,1,NA,36.869584,-118.189241,0,20.25,0,0,None,734,0,0,0,0,10,0,0.0,131.6,0.0,202.5,1,0,93526
754,0,0,1,0,2,1,0,Fiber optic,1,1,1,0,Month-to-month,0,Electronic check,90.35,190.5,0,19,53,4.65,5361,0,Temecula,0,0,Fiber Optic,33.507255,-117.029473,1,90.35,0,10,None,46171,0,0,1,0,2,2,101.0,9.3,0.0,190.5,1,0,92592
755,1,1,0,0,20,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.55,1842.8,1,73,14,44.44,5444,1,San Diego,1,1,Cable,32.961064,-117.13491699999999,0,102.492,0,0,None,47224,0,0,0,0,20,5,258.0,888.8,0.0,1842.8,0,0,92129
756,1,0,0,0,66,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.7,1253.8,0,50,0,45.54,4601,0,June Lake,0,1,NA,37.730269,-119.05581299999999,0,19.7,0,0,Offer A,618,0,0,0,0,66,2,0.0,3005.64,0.0,1253.8,0,0,93529
757,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,57.2,0,22,0,3.12,5634,0,Keeler,0,0,NA,36.560497999999995,-117.962461,0,19.85,0,0,None,71,0,0,0,0,3,0,0.0,9.36,0.0,57.2,1,0,93530
758,0,0,0,1,15,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),85.9,1269.55,1,37,14,24.63,3579,1,Keene,0,0,Cable,35.214982,-118.59048999999999,0,89.33600000000001,0,0,None,1436,0,0,0,1,15,2,178.0,369.45,0.0,1269.55,0,0,93531
759,0,0,1,1,72,1,1,Fiber optic,1,1,0,0,Two year,1,Bank transfer (automatic),90.35,6563.4,0,41,25,9.6,5794,0,Lake Hughes,0,0,Fiber Optic,34.659579,-118.58421200000001,1,90.35,0,9,Offer A,2771,1,0,1,0,72,1,0.0,691.1999999999998,0.0,6563.4,0,1,93532
760,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.8,20.8,0,37,0,48.14,3678,0,Lancaster,0,1,NA,34.727529,-118.153098,0,20.8,0,0,Offer E,35109,0,1,0,0,1,2,0.0,48.14,0.0,20.8,0,0,93534
761,0,0,0,0,22,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,89.25,1907.85,1,38,2,18.01,3161,1,Lancaster,0,0,Cable,34.712708,-117.889656,0,92.82,0,0,None,57794,0,2,0,1,22,2,0.0,396.22,0.0,1907.85,0,1,93535
762,1,0,1,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,208.85,1,31,12,26.71,3038,1,Lancaster,0,1,Cable,34.741406,-118.38111,1,73.112,0,1,None,49309,0,4,1,0,3,1,25.0,80.13,0.0,208.85,0,0,93536
763,0,0,1,1,72,1,1,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),66.85,4758.8,0,56,20,14.65,6264,0,Lee Vining,1,0,Fiber Optic,37.890145000000004,-119.184087,1,66.85,0,6,Offer A,504,1,0,1,0,72,3,952.0,1054.8,0.0,4758.8,0,0,93541
764,1,0,1,1,65,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.9,1292.6,0,30,0,18.07,6312,0,Littlerock,0,1,NA,34.505272999999995,-117.955054,1,19.9,0,2,Offer B,11198,0,0,1,0,65,1,0.0,1174.55,0.0,1292.6,0,0,93543
765,0,0,0,0,11,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Mailed check,35.8,363.15,0,22,52,0.0,2534,0,Llano,0,0,Fiber Optic,34.500091,-117.76586200000001,0,35.8,0,0,Offer D,1220,0,0,0,0,11,1,0.0,0.0,0.0,363.15,1,1,93544
766,1,0,0,0,22,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,78.85,1600.25,0,56,10,30.35,2444,0,Fallbrook,0,1,Cable,33.362575,-117.299644,0,78.85,0,0,Offer D,42239,0,0,0,0,22,2,160.0,667.7,0.0,1600.25,0,0,92028
767,1,0,0,0,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.4,275.7,0,23,0,36.42,5068,0,Mammoth Lakes,0,1,NA,37.550074,-118.837167,0,20.4,0,0,Offer D,8217,0,0,0,0,14,0,0.0,509.88,0.0,275.7,1,0,93546
768,1,0,0,0,41,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.25,3089.1,0,45,6,1.08,3277,0,Olancha,0,1,Fiber Optic,36.296851000000004,-117.86546899999999,0,74.25,0,0,Offer B,318,1,0,0,0,41,0,0.0,44.28,0.0,3089.1,0,1,93549
769,1,0,1,0,17,1,0,DSL,1,1,0,1,One year,0,Mailed check,64.8,1175.6,0,32,11,45.35,3546,0,Palmdale,0,1,Fiber Optic,34.536232,-118.082935,1,64.8,0,2,Offer D,67232,0,0,1,1,17,0,129.0,770.95,0.0,1175.6,0,0,93550
770,1,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.45,237.3,0,63,0,44.53,2642,0,Palmdale,0,1,NA,34.613476,-118.256358,0,20.45,0,0,Offer D,34045,0,0,0,0,11,0,0.0,489.83,0.0,237.3,0,0,93551
771,1,0,0,0,15,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.35,1444.65,1,49,16,48.93,5264,1,Palmdale,0,1,Cable,34.557711,-118.02944099999999,0,97.084,0,0,None,25370,0,1,0,1,15,1,231.0,733.95,0.0,1444.65,0,0,93552
772,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,19.9,1,45,0,49.51,4248,1,Pearblossom,0,0,NA,34.445239,-117.89486799999999,0,19.9,0,0,None,1613,0,0,0,0,1,2,0.0,49.51,0.0,19.9,0,0,93553
773,0,0,1,0,5,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Mailed check,88.9,454.15,1,37,30,41.57,4356,1,Randsburg,1,0,DSL,35.405722,-117.773354,1,92.456,0,1,None,117,0,0,1,1,5,0,136.0,207.85,0.0,454.15,0,0,93554
774,1,0,1,0,33,1,0,Fiber optic,0,0,1,1,One year,1,Electronic check,95.8,3036.75,1,24,45,41.8,4161,1,Temecula,1,1,DSL,33.507255,-117.029473,1,99.632,0,1,Offer C,46171,0,0,1,1,33,0,1367.0,1379.4,0.0,3036.75,1,0,92592
775,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),110.65,8065.65,0,24,73,41.21,4259,0,Rosamond,1,0,Fiber Optic,34.903052,-118.41125100000001,1,110.65,0,5,Offer A,14931,0,0,1,1,72,0,0.0,2967.12,0.0,8065.65,1,1,93560
776,0,0,1,1,3,0,No phone service,DSL,0,1,0,1,Month-to-month,0,Mailed check,40.3,92.5,0,59,53,0.0,5651,0,Tehachapi,0,0,Fiber Optic,35.073777,-118.65211200000002,1,40.3,3,6,Offer E,25805,0,0,1,1,3,0,0.0,0.0,0.0,92.5,0,1,93561
777,1,0,0,0,2,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,82.0,184.65,1,42,15,41.18,3051,1,Temecula,0,1,Cable,33.507255,-117.029473,0,85.28,0,0,None,46171,0,0,0,0,2,6,0.0,82.36,0.0,184.65,0,1,92592
778,0,0,1,0,59,1,1,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),107.0,6152.3,0,20,48,41.15,4620,0,Valyermo,1,0,DSL,34.39583,-117.734568,1,107.0,0,7,Offer B,413,1,0,1,1,59,1,2953.0,2427.85,0.0,6152.3,1,0,93563
779,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.35,89.5,1,63,10,25.49,3478,1,Palmdale,0,1,Cable,34.598221,-117.79593,0,47.163999999999994,0,0,None,6787,0,1,0,0,2,3,9.0,50.98,0.0,89.5,0,0,93591
780,1,0,1,1,71,1,0,DSL,0,1,1,1,Two year,1,Credit card (automatic),73.35,5154.5,0,30,59,16.24,5124,0,Ahwahnee,0,1,DSL,37.375816,-119.739935,1,73.35,0,4,Offer A,1968,1,0,1,1,71,0,0.0,1153.04,0.0,5154.5,0,1,93601
781,0,0,1,1,5,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.8,220.45,0,45,19,35.6,2492,0,Auberry,0,0,Fiber Optic,36.991762,-119.242874,1,44.8,2,10,Offer E,3464,0,0,1,0,5,1,0.0,178.0,0.0,220.45,0,1,93602
782,1,0,1,1,27,1,0,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),54.75,1510.3,0,54,53,36.19,3519,0,Badger,0,1,Fiber Optic,36.64545,-118.924982,1,54.75,6,5,None,273,0,0,1,0,27,2,800.0,977.13,0.0,1510.3,0,0,93603
783,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,52.2,52.2,1,41,25,34.04,4138,1,Bass Lake,0,0,Cable,37.458366999999996,-119.34501100000001,0,54.288,0,0,None,613,1,1,0,0,1,3,0.0,34.04,0.0,52.2,0,1,93604
784,1,0,0,1,63,0,No phone service,DSL,1,1,0,0,One year,1,Bank transfer (automatic),40.6,2588.95,0,48,28,0.0,6406,0,Big Creek,0,1,Fiber Optic,37.17277,-119.2997,0,40.6,0,0,Offer B,273,1,0,0,0,63,0,725.0,0.0,0.0,2588.95,0,0,93605
785,0,1,0,0,46,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,110.0,4874.8,1,65,22,2.37,2403,1,Biola,1,0,DSL,36.798882,-120.01951100000001,0,114.4,0,0,None,807,0,0,0,1,46,4,1072.0,109.02,0.0,4874.8,0,0,93606
786,1,0,1,1,72,1,1,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),55.3,3983.6,0,40,27,24.24,6259,0,Cantua Creek,0,1,DSL,36.488056,-120.40769099999999,1,55.3,0,5,Offer A,1766,0,0,1,0,72,1,0.0,1745.28,0.0,3983.6,0,1,93608
787,0,0,1,0,34,1,1,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),60.85,2003.6,0,59,26,12.3,3012,0,Caruthers,0,0,Cable,36.5276,-119.865999,1,60.85,0,5,None,5446,1,0,1,0,34,0,0.0,418.2000000000001,0.0,2003.6,0,1,93609
788,0,0,1,1,24,1,1,DSL,1,1,1,1,One year,0,Electronic check,78.4,1832.4,0,54,12,31.62,2506,0,Chowchilla,0,0,Fiber Optic,37.100947999999995,-120.27013600000001,1,78.4,0,4,None,19391,0,1,1,1,24,2,220.0,758.88,0.0,1832.4,0,0,93610
789,1,0,0,0,72,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),69.65,4908.25,0,53,13,3.66,4262,0,Clovis,1,1,Fiber Optic,36.917652000000004,-119.59375700000001,0,69.65,0,0,Offer A,46858,1,0,0,0,72,0,638.0,263.52,0.0,4908.25,0,0,93611
790,0,0,1,1,60,0,No phone service,DSL,1,0,1,1,Two year,0,Credit card (automatic),59.85,3590.2,0,46,19,0.0,5790,0,Clovis,1,0,Cable,36.814539,-119.711868,1,59.85,0,1,Offer B,33856,1,0,1,1,60,2,0.0,0.0,0.0,3590.2,0,1,93612
791,1,0,0,0,68,1,1,DSL,1,1,0,1,One year,1,Credit card (automatic),76.9,5023,0,60,13,1.27,5355,0,Coarsegold,1,1,Fiber Optic,37.212191,-119.749323,0,76.9,0,0,Offer A,9395,0,1,0,1,68,1,0.0,86.36,0.0,5023.0,0,1,93614
792,0,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.85,146.6,0,44,0,17.09,3260,0,Cutler,0,0,NA,36.497895,-119.28548400000001,1,19.85,0,8,Offer E,5519,0,0,1,0,8,0,0.0,136.72,0.0,146.6,0,0,93615
793,0,0,0,1,34,1,0,DSL,1,0,1,0,Two year,0,Credit card (automatic),67.65,2339.3,0,22,27,20.75,4263,0,Del Rey,1,0,Fiber Optic,36.657462,-119.595293,0,67.65,0,0,None,1965,1,0,0,0,34,0,0.0,705.5,0.0,2339.3,1,1,93616
794,0,0,0,0,6,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Credit card (automatic),45.0,298.7,0,25,52,0.0,2270,0,Dinuba,0,0,DSL,36.523619000000004,-119.38686799999999,0,45.0,0,0,Offer E,24206,0,0,0,1,6,0,155.0,0.0,0.0,298.7,1,0,93618
795,1,0,1,0,2,1,0,DSL,0,1,0,1,Month-to-month,1,Mailed check,64.2,143.65,0,38,26,4.41,4369,0,Dos Palos,0,1,Fiber Optic,37.045728000000004,-120.63068200000001,1,64.2,0,2,Offer E,9388,1,0,1,1,2,1,37.0,8.82,0.0,143.65,0,0,93620
796,1,0,0,0,31,1,1,Fiber optic,0,0,0,0,One year,0,Credit card (automatic),81.7,2548.65,0,24,76,17.18,4850,0,Dunlap,0,1,DSL,36.789213000000004,-119.14033799999999,0,81.7,0,0,None,506,1,0,0,0,31,0,1937.0,532.58,0.0,2548.65,1,0,93621
797,0,0,1,1,20,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),25.55,507.4,0,47,0,36.85,3235,0,Firebaugh,0,0,NA,36.785618,-120.625382,1,25.55,7,6,Offer D,9491,0,1,1,0,20,2,0.0,737.0,0.0,507.4,0,0,93622
798,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.0,20,0,21,0,6.86,2358,0,Fish Camp,0,0,NA,37.483534999999996,-119.679414,1,20.0,3,4,None,77,0,1,1,0,1,2,0.0,6.86,0.0,20.0,1,0,93623
799,1,0,0,0,62,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,96.75,6125.4,1,58,10,22.64,5016,1,Five Points,1,1,DSL,36.397745,-120.11991100000002,0,100.62,0,0,Offer B,1852,0,0,0,1,62,2,613.0,1403.68,0.0,6125.4,0,0,93624
800,0,1,1,0,70,1,1,Fiber optic,0,0,0,0,Two year,1,Credit card (automatic),75.65,5411.4,0,72,3,16.87,4181,0,Fowler,0,0,Fiber Optic,36.625792,-119.67248300000001,1,75.65,0,4,Offer A,5635,0,0,1,0,70,0,162.0,1180.9,25.67,5411.4,0,0,93625
801,0,0,0,0,10,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.5,1058.25,1,33,33,14.53,5184,1,Friant,0,0,Cable,37.027663000000004,-119.69056,0,102.44,0,0,None,1125,1,1,0,1,10,2,349.0,145.29999999999995,0.0,1058.25,0,0,93626
802,1,0,1,1,39,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,23.8,903.8,0,39,0,29.56,3970,0,Helm,0,1,NA,36.520537,-120.118055,1,23.8,0,7,None,152,0,0,1,0,39,0,0.0,1152.84,0.0,903.8,0,0,93627
803,0,0,1,0,46,1,0,DSL,0,1,1,0,Two year,1,Credit card (automatic),64.2,3009.5,0,61,6,37.02,4699,0,Hume,0,0,DSL,36.807595,-118.901544,1,64.2,0,1,None,93,1,0,1,0,46,3,0.0,1702.92,0.0,3009.5,0,1,93628
804,1,0,0,0,6,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,85.35,489.45,1,61,30,11.97,4694,1,Kerman,0,1,Cable,36.727418,-120.123526,0,88.764,0,0,None,14062,0,0,0,0,6,4,0.0,71.82000000000002,0.0,489.45,0,1,93630
805,0,0,1,1,72,1,1,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),76.8,5468.45,0,45,9,43.47,5120,0,Kingsburg,1,0,Fiber Optic,36.478239,-119.52136999999999,1,76.8,0,5,Offer A,14088,0,0,1,1,72,1,0.0,3129.84,0.0,5468.45,0,1,93631
806,1,0,0,0,18,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),55.2,1058.1,0,63,28,47.72,2110,0,Lakeshore,1,1,Fiber Optic,37.290606,-119.216328,0,55.2,0,0,Offer D,52,1,0,0,0,18,0,0.0,858.96,0.0,1058.1,0,1,93634
807,1,0,1,0,71,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),108.55,7616,0,29,73,31.97,4111,0,Los Banos,1,1,Fiber Optic,36.995162,-120.955099,1,108.55,0,10,Offer A,29124,1,0,1,1,71,0,0.0,2269.87,0.0,7616.0,1,1,93635
808,1,0,1,0,40,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.3,4113.1,1,54,4,22.56,2576,1,Madera,0,1,Fiber Optic,36.902954,-120.194274,1,105.352,0,1,Offer B,28434,0,3,1,1,40,4,0.0,902.4,0.0,4113.1,0,1,93637
809,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.55,69.55,1,27,53,49.43,3042,1,Madera,0,1,DSL,37.004068,-119.930027,0,72.332,0,0,Offer E,49247,0,0,0,1,1,7,0.0,49.43,0.0,69.55,1,0,93638
810,1,0,0,0,58,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),103.25,6017.65,1,20,52,44.5,6105,1,Escondido,1,1,Cable,33.141265000000004,-116.967221,0,107.38,0,0,Offer B,48690,0,1,0,1,58,1,0.0,2581.0,0.0,6017.65,1,1,92027
811,1,0,0,0,70,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),104.0,7250.15,1,25,46,12.19,4544,1,Miramonte,0,1,DSL,36.696759,-119.024051,0,108.16,0,0,Offer A,571,1,0,0,1,70,5,3335.0,853.3,0.0,7250.15,1,0,93641
812,0,0,1,0,42,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,25.25,1108.2,0,55,0,33.63,3052,0,North Fork,0,0,NA,37.244307,-119.470256,1,25.25,0,9,None,3376,0,0,1,0,42,1,0.0,1412.46,0.0,1108.2,0,0,93643
813,1,0,1,1,34,0,No phone service,DSL,1,0,0,0,One year,0,Bank transfer (automatic),30.4,938.65,0,23,42,0.0,4697,0,Oakhurst,0,1,Cable,37.648647,-119.231447,1,30.4,0,0,None,8521,0,0,0,0,34,0,0.0,0.0,0.0,938.65,1,1,93644
814,1,1,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.05,94.15,0,65,0,30.14,2154,0,O Neals,0,1,NA,37.140104,-119.65709199999999,0,20.05,0,0,Offer E,173,0,0,0,0,5,0,0.0,150.7,0.0,94.15,0,0,93645
815,0,0,0,0,25,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,84.6,2088.05,0,23,59,9.57,4874,0,Orange Cove,0,0,DSL,36.633497999999996,-119.298895,0,84.6,0,0,Offer C,8449,0,0,0,0,25,0,1232.0,239.25,0.0,2088.05,1,0,93646
816,0,0,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Mailed check,86.2,178.7,1,62,30,24.05,2969,1,Orosi,1,0,Cable,36.600184999999996,-119.175655,0,89.64800000000002,0,0,Offer E,9780,0,0,0,1,2,2,0.0,48.1,0.0,178.7,0,1,93647
817,0,0,1,1,55,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),103.7,5656.75,0,37,57,35.04,5892,0,Parlier,1,0,Cable,36.622237,-119.521126,1,103.7,3,10,None,12587,1,0,1,1,55,0,0.0,1927.2,0.0,5656.75,0,1,93648
818,1,0,1,0,21,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,111.2,2317.1,1,24,65,36.26,4123,1,Fresno,1,1,Fiber Optic,36.841654999999996,-119.79711299999998,1,115.648,0,1,None,3258,1,0,1,1,21,1,150.61,761.4599999999998,0.0,2317.1,1,1,93650
819,1,0,1,0,70,1,1,Fiber optic,1,1,0,0,Two year,1,Credit card (automatic),88.0,5986.45,0,30,51,9.28,4867,0,Prather,0,1,DSL,37.007238,-119.505661,1,88.0,0,9,None,1314,1,0,1,0,70,2,3053.0,649.5999999999998,0.0,5986.45,0,0,93651
820,0,0,1,0,61,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,106.35,6751.35,0,41,29,27.63,5632,0,Raisin City,1,0,Fiber Optic,36.594542,-119.905245,1,106.35,0,3,None,265,1,0,1,1,61,0,0.0,1685.4299999999996,0.0,6751.35,0,1,93652
821,1,0,1,1,43,1,0,DSL,1,0,1,1,Two year,1,Credit card (automatic),79.15,3566.6,0,62,18,41.08,3716,0,Raymond,1,1,Cable,37.252057,-119.95783,1,79.15,0,1,None,972,1,0,1,1,43,2,642.0,1766.4399999999996,0.0,3566.6,0,0,93653
822,1,0,0,0,47,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,103.1,4889.3,0,37,8,16.64,5029,0,Reedley,1,1,Cable,36.636638,-119.421842,0,103.1,0,0,None,25923,0,1,0,1,47,3,391.0,782.08,0.0,4889.3,0,0,93654
823,1,0,0,0,5,1,0,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),63.95,318.1,0,38,5,13.96,3099,0,Riverdale,1,1,Fiber Optic,36.452211,-119.94575,0,63.95,0,0,Offer E,5729,1,0,0,0,5,0,0.0,69.80000000000001,0.0,318.1,0,1,93656
824,0,0,0,0,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.8,1563.95,0,55,0,8.23,6201,0,Sanger,0,0,NA,36.819628,-119.44041399999999,0,25.8,0,0,None,28991,0,0,0,0,62,1,0.0,510.2600000000001,0.0,1563.95,0,0,93657
825,0,0,1,1,16,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),89.45,1430.25,1,41,28,31.73,3696,1,San Joaquin,1,0,DSL,36.600193,-120.153393,1,93.02799999999999,0,1,None,4318,0,0,1,0,16,2,400.0,507.68,0.0,1430.25,0,0,93660
826,1,1,1,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.6,644.35,1,74,12,21.91,3265,1,Selma,0,1,Cable,36.545322,-119.64228100000001,1,99.424,0,1,None,26213,0,0,1,0,7,1,77.0,153.37,0.0,644.35,0,0,93662
827,0,0,1,1,14,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,25.55,372.45,0,47,0,31.7,2080,0,Shaver Lake,0,0,NA,37.223,-119.001021,1,25.55,1,1,None,642,0,0,1,0,14,2,0.0,443.8,0.0,372.45,0,0,93664
828,1,0,1,1,60,1,0,Fiber optic,0,1,1,0,One year,0,Electronic check,90.95,5453.4,1,21,57,33.25,4111,1,South Dos Palos,1,1,Cable,36.959731,-120.65351899999999,1,94.588,0,1,Offer B,343,0,0,1,1,60,3,0.0,1995.0,0.0,5453.4,1,1,93665
829,1,0,1,1,34,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,44.85,1442.6,0,35,76,0.0,5569,0,Sultana,1,1,Fiber Optic,36.545353000000006,-119.33853500000001,1,44.85,3,2,Offer C,306,1,0,1,0,34,1,0.0,0.0,0.0,1442.6,0,1,93666
830,0,0,1,0,50,1,1,Fiber optic,1,1,1,1,One year,0,Electronic check,108.55,5610.7,1,58,15,29.43,4274,1,Tollhouse,0,0,Cable,36.993666,-119.34826699999999,1,112.89200000000001,0,1,Offer B,2633,1,0,1,1,50,3,842.0,1471.5,0.0,5610.7,0,0,93667
831,1,0,1,1,38,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.05,963.95,0,44,0,33.1,3772,0,Tranquillity,0,1,NA,36.635661,-120.28864399999999,1,25.05,1,9,Offer C,1130,0,0,1,0,38,2,0.0,1257.8,0.0,963.95,0,0,93668
832,0,0,1,1,70,1,0,DSL,1,1,0,1,One year,0,Credit card (automatic),74.1,5222.3,0,46,21,19.1,6325,0,Wishon,1,0,Fiber Optic,37.287758000000004,-119.548156,1,74.1,0,7,None,327,1,0,1,1,70,0,1097.0,1337.0,0.0,5222.3,0,0,93669
833,0,0,1,1,37,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,88.8,3340.55,0,33,16,1.08,3746,0,Traver,0,0,Fiber Optic,36.456091,-119.486225,1,88.8,2,3,Offer C,646,0,0,1,0,37,1,534.0,39.96,0.0,3340.55,0,0,93673
834,0,1,0,0,4,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,78.85,292.8,1,65,20,36.93,5301,1,Squaw Valley,0,0,Cable,36.719141,-119.20267700000001,0,82.00399999999998,0,0,None,3146,0,2,0,0,4,3,59.0,147.72,0.0,292.8,0,0,93675
835,1,1,1,1,60,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,93.25,5774.55,0,70,53,19.68,4353,0,Fresno,0,1,Fiber Optic,36.749403,-119.78757399999999,1,93.25,3,4,None,13858,0,0,1,0,60,1,0.0,1180.8,0.0,5774.55,0,1,93701
836,1,0,1,1,62,1,0,DSL,1,0,0,1,One year,0,Credit card (automatic),71.4,4487.3,0,47,25,14.05,5327,0,Fresno,1,1,Fiber Optic,36.739385,-119.753649,1,71.4,0,0,None,47999,1,0,0,1,62,0,0.0,871.1,0.0,4487.3,0,1,93702
837,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.4,44.4,1,45,13,32.44,3522,1,Fresno,0,1,DSL,36.768774,-119.76263300000001,0,46.176,0,0,Offer E,31180,0,2,0,0,1,2,0.0,32.44,0.0,44.4,0,0,93703
838,1,0,0,0,36,1,0,DSL,1,0,1,1,Month-to-month,1,Credit card (automatic),79.2,2854.95,0,27,52,42.51,4830,0,Fresno,1,1,DSL,36.799648,-119.801247,0,79.2,0,0,Offer C,26580,1,0,0,1,36,0,1485.0,1530.36,0.0,2854.95,1,0,93704
839,1,0,0,0,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.4,905.55,0,36,0,1.4,2404,0,Fresno,0,1,NA,36.787240000000004,-119.82781299999999,0,20.4,0,0,None,35451,0,0,0,0,44,0,0.0,61.6,0.0,905.55,0,0,93705
840,0,1,0,0,55,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,100.0,5509.3,1,66,8,37.38,5679,1,Fresno,1,0,Cable,36.654614,-119.903674,0,104.0,0,0,None,35790,0,0,0,1,55,6,441.0,2055.9,0.0,5509.3,0,0,93706
841,0,0,1,0,72,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),105.0,7589.8,0,44,7,6.58,5678,0,Fresno,1,0,DSL,36.822715,-119.761826,1,105.0,0,7,None,29337,0,0,1,1,72,1,0.0,473.76,0.0,7589.8,0,1,93710
842,0,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.8,229.6,1,59,0,37.65,2653,1,Fresno,0,0,NA,36.833002,-119.82947,1,19.8,0,1,None,36274,0,0,1,0,12,4,0.0,451.8,0.0,229.6,0,0,93711
843,0,0,0,0,13,0,No phone service,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),30.85,394.1,0,59,7,0.0,2444,0,Fresno,0,0,Fiber Optic,36.878709,-119.7645,0,30.85,0,0,None,45087,0,0,0,0,13,0,28.0,0.0,0.0,394.1,0,0,93720
844,1,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.9,89.9,1,21,58,32.85,5951,1,Fresno,0,1,Cable,36.732694,-119.783786,0,93.496,0,0,Offer E,6848,0,0,0,1,1,1,0.0,32.85,0.0,89.9,1,0,93721
845,0,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.55,295.95,0,23,0,34.63,3009,0,Fresno,0,0,NA,36.78979,-119.92989399999999,1,20.55,0,7,None,60889,0,0,1,0,15,1,0.0,519.45,0.0,295.95,1,0,93722
846,0,0,0,0,65,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),84.85,5459.2,0,57,17,41.74,5434,0,Fresno,1,0,DSL,36.623632,-119.741322,0,84.85,0,0,None,21010,1,0,0,1,65,0,0.0,2713.1,0.0,5459.2,0,1,93725
847,0,0,1,1,12,0,No phone service,DSL,1,0,0,0,One year,0,Credit card (automatic),33.15,444.75,0,54,27,0.0,3882,0,Fresno,0,0,DSL,36.793601,-119.761131,1,33.15,0,7,None,39148,1,0,1,0,12,1,0.0,0.0,0.0,444.75,0,1,93726
848,1,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),92.0,6782.15,0,55,5,5.32,5883,0,Fresno,1,1,Fiber Optic,36.751489,-119.68072,1,92.0,0,8,None,54701,1,0,1,1,72,3,0.0,383.04,0.0,6782.15,0,1,93727
849,0,0,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.8,6510.45,0,23,69,44.92,5762,0,Fresno,1,0,DSL,36.757345,-119.818274,1,89.8,0,3,None,16346,1,0,1,1,72,1,4492.0,3234.24,0.0,6510.45,1,0,93728
850,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),115.8,8476.5,0,57,24,12.29,5841,0,Salinas,1,0,Fiber Optic,36.64152,-121.622188,1,115.8,2,9,None,35739,1,0,1,1,72,0,0.0,884.8799999999999,0.0,8476.5,0,1,93901
851,1,0,0,1,52,1,1,DSL,1,1,1,1,Two year,1,Mailed check,85.15,4461.85,0,63,28,32.02,4322,0,Salinas,0,1,DSL,36.667794,-121.60130600000001,0,85.15,0,0,None,58548,1,1,0,1,52,3,124.93,1665.0400000000004,0.0,4461.85,0,1,93905
852,1,0,0,0,2,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,24.85,62,0,50,0,40.25,5983,0,Salinas,0,1,NA,36.722898,-121.633648,0,24.85,0,0,Offer E,53946,0,0,0,0,2,0,0.0,80.5,0.0,62.0,0,0,93906
853,0,0,0,0,5,1,0,DSL,1,0,1,0,Month-to-month,1,Electronic check,64.35,352.65,0,63,22,8.32,4771,0,Salinas,0,0,Fiber Optic,36.77462,-121.66471399999999,0,64.35,0,0,Offer E,22292,1,0,0,0,5,1,78.0,41.6,0.0,352.65,0,0,93907
854,0,0,0,0,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.5,1424.9,0,32,0,48.41,4201,0,Salinas,0,0,NA,36.624338,-121.615669,0,20.5,0,0,None,13027,0,0,0,0,68,2,0.0,3291.88,0.0,1424.9,0,0,93908
855,0,0,0,1,62,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,100.15,6413.65,1,41,16,32.58,5600,1,Escondido,1,0,Cable,33.141265000000004,-116.967221,0,104.156,0,0,Offer B,48690,0,0,0,1,62,5,1026.0,2019.96,0.0,6413.65,0,0,92027
856,1,0,0,0,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),86.05,6309.65,0,22,71,48.36,5965,0,Carmel By The Sea,0,1,DSL,36.554618,-121.92223899999999,0,86.05,0,0,None,2966,1,0,0,1,72,0,447.99,3481.92,0.0,6309.65,1,1,93921
857,1,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,50.8,50.8,1,58,30,1.28,3718,1,Carmel,0,1,DSL,36.460611,-121.852507,0,52.832,0,0,Offer E,13121,0,2,0,0,1,3,0.0,1.28,0.0,50.8,0,0,93923
858,0,0,1,0,66,1,1,Fiber optic,1,1,0,0,One year,0,Electronic check,89.0,5898.6,0,59,8,37.38,4488,0,Carmel Valley,0,0,Fiber Optic,36.414611,-121.6386,1,89.0,0,10,None,6691,1,0,1,0,66,0,0.0,2467.080000000001,0.0,5898.6,0,1,93924
859,1,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,1,Credit card (automatic),64.8,4719.75,0,52,18,0.0,4036,0,Chualar,1,1,DSL,36.596271,-121.442274,1,64.8,0,9,None,1140,1,0,1,1,72,0,850.0,0.0,0.0,4719.75,0,0,93925
860,1,0,0,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.8,457.3,0,63,0,45.7,5823,0,Gonzales,0,1,NA,36.52588,-121.39671899999999,0,19.8,0,0,Offer C,9023,0,1,0,0,26,2,0.0,1188.2,0.0,457.3,0,0,93926
861,1,0,1,1,64,1,1,Fiber optic,1,0,0,1,Two year,0,Bank transfer (automatic),93.4,5822.3,0,53,11,30.82,6249,0,Greenfield,1,1,Fiber Optic,36.248708,-121.38661699999999,1,93.4,1,2,None,14204,0,0,1,1,64,1,640.0,1972.48,0.0,5822.3,0,0,93927
862,1,1,1,0,20,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,73.65,1463.5,1,71,26,5.37,5849,1,Jolon,0,1,Cable,35.930782,-121.189757,1,76.596,0,1,None,254,0,0,1,0,20,0,0.0,107.4,0.0,1463.5,0,1,93928
863,0,0,0,0,3,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,95.1,307.4,1,55,32,47.62,5861,1,King City,0,0,Fiber Optic,36.220760999999996,-120.980777,0,98.904,0,0,Offer E,14477,0,1,0,1,3,2,0.0,142.86,0.0,307.4,0,1,93930
864,1,0,0,0,22,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),94.65,2104.55,1,52,18,46.28,3665,1,Lockwood,0,1,DSL,35.989792,-121.05593300000001,0,98.436,0,0,None,538,0,0,0,1,22,4,379.0,1018.16,0.0,2104.55,0,0,93932
865,1,0,1,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,80.6,319.15,1,46,2,14.3,3080,1,Marina,1,1,Cable,36.689582,-121.758398,1,83.824,0,1,Offer E,21759,1,0,1,0,4,0,6.0,57.2,0.0,319.15,0,0,93933
866,1,0,1,0,62,0,No phone service,DSL,0,0,1,0,Two year,1,Bank transfer (automatic),39.0,2337.45,0,61,4,0.0,4987,0,Monterey,0,1,Cable,36.362741,-121.869685,1,39.0,0,6,None,32857,1,0,1,0,62,2,93.0,0.0,0.0,2337.45,0,0,93940
867,0,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.5,104.3,0,44,0,24.61,5263,0,Pacific Grove,0,0,NA,36.618337,-121.92641699999999,0,20.5,0,0,None,15449,0,0,0,0,5,0,0.0,123.05,0.0,104.3,0,0,93950
868,1,0,1,0,59,1,1,Fiber optic,0,0,0,1,One year,0,Electronic check,85.55,5084.65,1,24,57,6.91,6304,1,Pebble Beach,0,1,Fiber Optic,36.587497,-121.94481499999999,1,88.97200000000001,0,0,Offer B,4602,0,1,0,1,59,4,2898.0,407.69,0.0,5084.65,1,0,93953
869,1,0,0,1,3,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,26.4,121.25,0,44,0,33.87,4315,0,San Lucas,0,1,NA,36.125529,-120.864443,0,26.4,1,0,None,521,0,0,0,0,3,0,0.0,101.61,0.0,121.25,0,0,93954
870,0,0,1,0,72,1,1,Fiber optic,1,0,1,0,Two year,1,Bank transfer (automatic),98.2,7015.9,0,32,3,25.48,4332,0,Seaside,1,0,Fiber Optic,36.625114,-121.82356499999999,1,98.2,0,1,None,38244,1,0,1,0,72,1,210.0,1834.56,0.0,7015.9,0,0,93955
871,1,0,1,1,57,1,0,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),97.55,5598,0,26,73,4.18,5833,0,Soledad,1,1,DSL,36.414215999999996,-121.360597,1,97.55,3,1,None,13003,0,0,1,1,57,1,4087.0,238.26,0.0,5598.0,1,0,93960
872,1,0,0,1,66,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.95,1269.1,0,63,0,37.94,6382,0,Spreckels,0,1,NA,36.624641,-121.647195,0,19.95,1,0,None,407,0,0,0,0,66,2,0.0,2504.04,0.0,1269.1,0,0,93962
873,0,0,0,0,60,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,50.8,3027.4,1,58,6,0.0,4941,1,Belmont,0,0,DSL,37.509366,-122.306132,0,52.832,0,0,Offer B,25566,0,0,0,1,60,0,182.0,0.0,0.0,3027.4,0,0,94002
874,1,0,0,1,45,1,1,Fiber optic,0,0,1,1,Two year,0,Bank transfer (automatic),99.7,4634.35,0,33,12,23.54,3333,0,Brisbane,1,1,Fiber Optic,37.684694,-122.40711999999999,0,99.7,2,0,None,3635,0,0,0,1,45,0,0.0,1059.3,0.0,4634.35,0,1,94005
875,0,0,0,0,3,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),34.8,113.95,0,25,46,0.0,2496,0,Burlingame,0,0,Cable,37.57028,-122.365778,0,34.8,0,0,None,40346,0,0,0,0,3,0,0.0,0.0,0.0,113.95,1,1,94010
876,0,0,0,0,15,1,0,Fiber optic,1,0,1,1,Month-to-month,0,Electronic check,105.1,1582.75,1,54,8,22.39,2122,1,Daly City,1,0,DSL,37.691561,-122.445202,0,109.304,0,0,None,47453,1,0,0,1,15,5,127.0,335.85,0.0,1582.75,0,0,94014
877,0,0,0,1,51,0,No phone service,DSL,1,0,1,1,One year,0,Bank transfer (automatic),60.15,3077,0,48,10,0.0,5404,0,Daly City,1,0,Cable,37.680844,-122.48131000000001,0,60.15,0,0,None,63337,1,0,0,1,51,2,0.0,0.0,0.0,3077.0,0,1,94015
878,0,0,0,0,60,1,1,DSL,1,0,0,0,One year,0,Electronic check,64.75,4039.5,0,29,27,37.95,6408,0,Half Moon Bay,1,0,Fiber Optic,37.45567,-122.407992,0,64.75,0,0,None,17929,1,0,0,0,60,0,1091.0,2277.0,0.0,4039.5,1,0,94019
879,1,0,0,0,33,1,1,DSL,0,1,0,0,Month-to-month,1,Bank transfer (automatic),54.65,1665.2,0,62,5,5.91,5201,0,La Honda,0,1,DSL,37.285677,-122.22416499999999,0,54.65,0,0,Offer C,1622,0,1,0,0,33,1,0.0,195.03,0.0,1665.2,0,1,94020
880,1,0,0,0,10,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,110.1,1043.3,1,53,7,18.03,5803,1,Loma Mar,1,1,DSL,37.266388,-122.26308,0,114.50399999999999,0,0,None,148,1,1,0,1,10,5,7.3,180.3,0.0,1043.3,0,1,94021
881,1,1,0,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.3,504.2,0,65,0,29.88,2269,0,Los Altos,0,1,NA,37.349546000000004,-122.13435600000001,0,19.3,0,0,Offer C,18486,0,0,0,0,26,0,0.0,776.88,9.49,504.2,0,0,94022
882,0,0,0,0,6,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,83.9,497.55,1,40,26,25.93,3962,1,Los Altos,1,0,DSL,37.352911,-122.093002,0,87.25600000000001,0,0,None,21496,0,0,0,1,6,0,129.0,155.57999999999996,0.0,497.55,0,0,94024
883,0,0,1,0,67,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,111.25,7511.65,0,39,23,35.03,5649,0,Menlo Park,1,0,DSL,37.449551,-122.18376200000002,1,111.25,0,1,None,39062,1,0,1,1,67,1,0.0,2347.01,0.0,7511.65,0,1,94025
884,0,0,1,1,49,0,No phone service,DSL,1,0,0,0,One year,1,Credit card (automatic),35.8,1782,0,19,82,0.0,4865,0,Atherton,0,0,DSL,37.454924,-122.20316799999999,1,35.8,0,1,None,6876,1,0,1,0,49,0,0.0,0.0,0.0,1782.0,1,1,94027
885,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.05,20.05,0,42,0,3.23,5368,0,Portola Valley,0,1,NA,37.369709,-122.21584399999999,0,20.05,0,0,None,6601,0,0,0,0,1,2,0.0,3.23,0.0,20.05,0,0,94028
886,0,1,0,0,7,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.35,609.65,0,66,20,26.29,2107,0,Millbrae,1,0,Cable,37.601248,-122.403099,0,84.35,0,0,Offer E,20350,0,0,0,0,7,0,0.0,184.03,29.17,609.65,0,1,94030
887,0,1,0,0,27,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),110.5,2857.6,0,70,4,35.76,4997,0,Montara,1,0,DSL,37.540582,-122.50959399999999,0,110.5,0,0,Offer C,2346,0,0,0,0,27,0,114.0,965.52,0.0,2857.6,0,0,94037
888,1,0,1,1,37,1,0,Fiber optic,0,0,1,1,One year,0,Credit card (automatic),91.2,3247.55,0,23,51,43.01,5263,0,Moss Beach,0,1,Cable,37.515556,-122.502311,1,91.2,3,1,Offer C,3064,0,1,1,1,37,1,165.63,1591.37,0.0,3247.55,1,1,94038
889,0,0,1,1,63,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,100.55,6215.35,1,48,18,8.98,5413,1,Mountain View,1,0,DSL,37.380662,-122.086022,1,104.572,0,3,Offer B,32143,0,0,1,0,63,0,1119.0,565.74,0.0,6215.35,0,0,94040
890,1,0,1,1,31,1,1,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,89.3,2823,0,37,57,20.76,2132,0,Mountain View,1,1,Fiber Optic,37.388349,-122.075299,1,89.3,3,1,Offer C,13483,1,0,1,0,31,0,0.0,643.5600000000002,0.0,2823.0,0,1,94041
891,1,0,1,1,50,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),103.85,5017.9,1,55,15,42.21,5812,1,Mountain View,1,1,Fiber Optic,37.419725,-122.062947,1,108.004,0,6,Offer B,27822,0,0,1,1,50,6,753.0,2110.5,0.0,5017.9,0,0,94043
892,1,1,0,0,32,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),81.1,2619.25,0,77,5,1.12,2143,0,Pacifica,1,1,Cable,37.573633,-122.45516699999999,0,81.1,0,0,Offer C,38885,0,0,0,0,32,0,13.1,35.84,19.25,2619.25,0,1,94044
893,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,24.6,24.6,1,39,13,0.0,5768,1,Pescadero,0,0,Cable,37.22565,-122.297533,0,25.584000000000003,0,0,None,2055,0,0,0,0,1,1,0.0,0.0,0.0,24.6,0,0,94060
894,0,0,1,0,63,1,1,Fiber optic,0,0,0,0,One year,1,Credit card (automatic),81.2,4965.1,0,56,27,38.85,6063,0,Redwood City,0,0,Cable,37.461251000000004,-122.23541399999999,1,81.2,0,1,Offer B,35737,1,0,1,0,63,1,0.0,2447.55,0.0,4965.1,0,1,94061
895,1,0,0,0,30,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Credit card (automatic),94.3,2679.7,0,53,28,41.66,4219,0,Redwood City,0,1,Fiber Optic,37.410567,-122.297152,0,94.3,0,0,Offer C,25569,0,0,0,1,30,0,750.0,1249.8,0.0,2679.7,0,0,94062
896,1,0,1,0,71,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),116.1,8310.55,0,29,27,33.83,5027,0,Redwood City,1,1,DSL,37.499411,-122.19631799999999,1,116.1,0,1,None,32368,1,0,1,1,71,0,0.0,2401.93,0.0,8310.55,1,1,94063
897,0,0,0,0,53,1,1,Fiber optic,0,1,1,1,Two year,0,Electronic check,105.55,5682.25,0,33,19,12.92,5731,0,Redwood City,1,0,Fiber Optic,37.527497,-122.23094099999999,0,105.55,0,0,Offer B,10658,0,0,0,1,53,0,1080.0,684.76,0.0,5682.25,0,0,94065
898,0,0,0,0,12,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),98.9,1120.95,1,64,25,34.92,5559,1,San Bruno,0,0,Fiber Optic,37.624435999999996,-122.43066100000001,0,102.856,0,0,None,39566,1,1,0,1,12,5,28.02,419.04,0.0,1120.95,0,1,94066
899,1,0,1,0,50,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Credit card (automatic),94.4,4914.9,0,27,47,17.58,5548,0,San Carlos,0,1,DSL,37.497915,-122.26736100000001,1,94.4,0,1,Offer B,28098,0,0,1,1,50,3,0.0,878.9999999999999,0.0,4914.9,1,1,94070
900,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.5,27.55,0,19,0,27.17,4836,0,San Gregorio,0,0,NA,37.331762,-122.341444,0,19.5,0,0,None,291,0,0,0,0,2,0,0.0,54.34,0.0,27.55,1,0,94074
901,0,0,0,0,9,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Credit card (automatic),98.3,923.5,1,27,90,38.76,2954,1,South San Francisco,1,0,Cable,37.654436,-122.426468,0,102.23200000000001,0,0,None,60599,0,0,0,1,9,1,831.0,348.84,0.0,923.5,1,0,94080
902,1,0,0,0,17,1,0,Fiber optic,1,0,1,1,Month-to-month,0,Electronic check,93.85,1625.65,1,36,14,4.51,4940,1,Sunnyvale,0,1,Fiber Optic,37.378541,-122.02045600000001,0,97.604,0,0,None,64010,0,0,0,1,17,1,228.0,76.67,0.0,1625.65,0,0,94086
903,0,0,1,0,56,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),105.6,6068.65,0,35,13,34.1,4196,0,Sunnyvale,1,0,Fiber Optic,37.3511,-122.03731100000002,1,105.6,0,1,Offer B,50070,0,0,1,1,56,0,0.0,1909.6,0.0,6068.65,0,1,94087
904,1,0,1,1,67,1,0,DSL,1,1,1,1,Two year,0,Credit card (automatic),81.35,5398.6,0,60,18,45.25,4219,0,Sunnyvale,1,1,Cable,37.421633,-122.00961299999999,1,81.35,0,1,None,16985,0,0,1,1,67,1,0.0,3031.75,0.0,5398.6,0,1,94089
905,1,1,0,0,9,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.5,918.6,1,65,16,48.71,4038,1,San Francisco,1,1,Cable,37.7795,-122.419233,0,104.52,0,0,None,28998,0,1,0,1,9,4,147.0,438.39,0.0,918.6,0,0,94102
906,1,0,0,0,4,1,0,DSL,0,0,1,0,Month-to-month,1,Electronic check,56.4,234.85,0,38,30,20.76,5344,0,San Francisco,0,1,Fiber Optic,37.773146999999994,-122.41128700000002,0,56.4,0,0,None,23036,0,0,0,0,4,1,70.0,83.04,0.0,234.85,0,0,94103
907,1,0,0,0,19,1,0,DSL,0,1,0,1,One year,1,Bank transfer (automatic),65.35,1231.85,0,61,6,41.79,2051,0,San Francisco,0,1,Cable,37.791222,-122.40224099999999,0,65.35,0,0,None,384,1,0,0,1,19,0,74.0,794.01,0.0,1231.85,0,0,94104
908,0,0,0,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,170.9,0,26,0,45.87,5919,0,San Francisco,0,0,NA,37.789168,-122.395009,0,19.95,3,0,None,2066,0,0,0,0,8,0,0.0,366.96,0.0,170.9,1,0,94105
909,0,0,0,0,71,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,111.25,7984.15,0,29,53,41.92,4361,0,San Francisco,1,0,DSL,37.768881,-122.395521,0,111.25,0,0,None,17372,1,0,0,1,71,0,4232.0,2976.32,0.0,7984.15,1,0,94107
910,1,1,0,0,10,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,72.85,688.65,1,69,26,5.46,3189,1,San Francisco,0,1,DSL,37.791998,-122.408653,0,75.764,0,0,None,13723,0,4,0,0,10,5,179.0,54.6,0.0,688.65,0,0,94108
911,0,1,0,0,15,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Credit card (automatic),89.0,1288.3,0,72,21,1.67,4452,0,San Francisco,0,0,Fiber Optic,37.794487,-122.42227,0,89.0,0,0,None,56330,0,2,0,0,15,1,0.0,25.05,45.69,1288.3,0,1,94109
912,1,0,1,1,72,1,1,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),106.1,7848.5,0,40,26,11.67,6283,0,San Francisco,1,1,Cable,37.750021000000004,-122.415201,1,106.1,1,1,None,74641,0,0,1,1,72,0,0.0,840.24,0.0,7848.5,0,1,94110
913,1,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.05,267,0,42,0,16.59,4018,0,San Francisco,0,1,NA,37.801776000000004,-122.402293,0,20.05,0,0,None,3337,0,0,0,0,12,1,0.0,199.08,0.0,267.0,0,0,94111
914,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.2,1798.9,0,22,0,28.06,6499,0,San Francisco,0,1,NA,37.720498,-122.443119,1,25.2,2,1,None,73117,0,0,1,0,72,0,0.0,2020.32,0.0,1798.9,1,0,94112
915,1,1,1,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.55,73.55,1,75,7,36.92,4369,1,San Francisco,0,1,Cable,37.758084999999994,-122.43480100000001,1,76.492,0,0,None,30587,0,0,0,0,1,2,0.0,36.92,0.0,73.55,0,1,94114
916,0,1,0,0,23,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),75.4,1643.55,0,67,25,17.62,2491,0,San Francisco,0,0,DSL,37.786031,-122.437301,0,75.4,0,0,None,33122,0,0,0,0,23,1,0.0,405.2600000000001,0.0,1643.55,0,1,94115
917,1,0,0,0,72,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),65.55,4807.45,0,45,10,0.0,4266,0,San Francisco,1,1,DSL,37.744409999999995,-122.486764,0,65.55,0,0,None,42959,1,0,0,1,72,0,481.0,0.0,0.0,4807.45,0,0,94116
918,0,0,0,0,26,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,80.7,2193,0,37,22,20.64,4501,0,San Francisco,1,0,Fiber Optic,37.770533,-122.445121,0,80.7,0,0,Offer C,38756,0,1,0,0,26,2,0.0,536.64,0.0,2193.0,0,1,94117
919,0,0,0,0,21,1,0,Fiber optic,0,1,1,1,One year,1,Mailed check,104.55,2239.4,0,48,27,36.31,3471,0,San Francisco,1,0,DSL,37.781304,-122.461522,0,104.55,0,0,None,38955,1,0,0,1,21,0,605.0,762.51,0.0,2239.4,0,0,94118
920,1,0,1,0,60,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),24.15,1505.9,0,23,0,16.42,4501,0,San Francisco,0,1,NA,37.776718,-122.49578100000001,1,24.15,0,1,Offer B,42476,0,0,1,0,60,2,0.0,985.2,0.0,1505.9,1,0,94121
921,1,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.45,255.35,0,26,0,41.11,4883,0,San Francisco,0,1,NA,37.760412,-122.48496599999999,0,20.45,0,0,None,55504,0,0,0,0,12,1,0.0,493.32,0.0,255.35,1,0,94122
922,1,0,1,0,16,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.4,1189.4,0,25,46,25.83,5432,0,San Francisco,0,1,Fiber Optic,37.800253999999995,-122.436975,1,75.4,0,1,None,22920,0,0,1,0,16,1,54.71,413.28,0.0,1189.4,1,1,94123
923,0,0,1,0,63,1,1,DSL,1,1,1,1,One year,1,Credit card (automatic),79.7,4786.15,0,38,24,49.08,4010,0,San Francisco,0,0,Cable,37.731505,-122.38453200000001,1,79.7,0,1,Offer B,33177,0,1,1,1,63,2,1149.0,3092.04,0.0,4786.15,0,0,94124
924,0,1,0,0,22,1,0,Fiber optic,1,1,0,0,Month-to-month,0,Electronic check,81.7,1820.9,0,77,22,23.43,5602,0,San Francisco,0,0,DSL,37.736534999999996,-122.45732,0,81.7,0,0,None,20643,0,0,0,0,22,3,401.0,515.46,29.88,1820.9,0,0,94127
925,0,0,1,1,32,1,0,DSL,1,1,0,1,Month-to-month,0,Bank transfer (automatic),76.3,2404.15,0,54,19,32.43,5324,0,San Francisco,1,0,Cable,37.797526,-122.46453100000001,1,76.3,1,1,Offer C,2240,1,0,1,1,32,0,45.68,1037.76,0.0,2404.15,0,1,94129
926,0,1,0,0,3,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.4,205.05,1,75,12,41.9,3501,1,San Francisco,0,0,Cable,37.820894,-122.369725,0,82.57600000000002,0,0,None,1458,0,1,0,0,3,5,25.0,125.7,0.0,205.05,0,0,94130
927,0,0,0,0,13,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,81.15,952.3,1,37,4,3.84,4806,1,San Francisco,1,0,DSL,37.746699,-122.44283300000001,0,84.39600000000002,0,0,None,27906,0,3,0,0,13,2,38.0,49.92,0.0,952.3,0,0,94131
928,0,0,1,1,68,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),103.75,7039.45,0,32,53,16.09,4121,0,San Francisco,0,0,Fiber Optic,37.722302,-122.491129,1,103.75,3,6,None,26297,1,0,1,1,68,0,3731.0,1094.12,0.0,7039.45,0,0,94132
929,0,0,1,1,30,1,0,Fiber optic,0,0,0,1,One year,0,Electronic check,86.45,2538.05,0,53,58,48.43,2923,0,San Francisco,1,0,DSL,37.802071000000005,-122.411004,1,86.45,3,0,Offer C,26831,0,0,0,1,30,0,0.0,1452.9,0.0,2538.05,0,1,94133
930,0,0,0,0,16,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),75.1,1212.85,0,44,25,38.02,5176,0,San Francisco,0,0,Fiber Optic,37.721052,-122.413573,0,75.1,0,0,None,40137,0,0,0,0,16,1,30.32,608.32,0.0,1212.85,0,1,94134
931,1,0,0,0,33,1,0,Fiber optic,0,1,0,0,Two year,0,Bank transfer (automatic),80.6,2651.1,0,32,27,34.85,5542,0,Palo Alto,0,1,DSL,37.444314,-122.149996,0,80.6,0,0,Offer C,16198,1,0,0,0,33,0,0.0,1150.05,0.0,2651.1,0,1,94301
932,1,0,1,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.3,1304.8,0,54,0,2.61,4035,0,Palo Alto,0,1,NA,37.458090000000006,-122.115398,1,19.3,0,3,None,45499,0,0,1,0,72,2,0.0,187.92,0.0,1304.8,0,0,94303
933,0,1,0,0,4,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.6,360.1,1,68,19,6.68,2467,1,Palo Alto,0,0,DSL,37.386978000000006,-122.177746,0,87.984,0,0,None,1723,0,1,0,0,4,6,6.84,26.72,0.0,360.1,0,1,94304
934,0,0,0,0,12,0,No phone service,DSL,1,0,0,0,One year,1,Mailed check,33.6,435.45,0,58,19,0.0,2990,0,Stanford,0,0,DSL,37.424341999999996,-122.165641,0,33.6,0,0,None,13386,1,0,0,0,12,0,83.0,0.0,0.0,435.45,0,0,94305
935,0,1,1,0,4,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,83.25,308.05,0,73,14,14.34,5251,0,Palo Alto,0,0,DSL,37.416159,-122.13133700000002,1,83.25,0,10,None,24492,0,1,1,0,4,3,43.0,57.36,39.93,308.05,0,0,94306
936,0,0,1,1,0,1,0,DSL,1,1,1,1,Two year,0,Mailed check,80.85, ,0,40,5,31.09,2048,0,San Mateo,1,0,Cable,37.590421,-122.306467,1,80.85,0,8,None,32488,0,0,1,1,10,2,40.0,310.9,0.0,808.5,0,0,94401
937,0,0,0,0,6,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,79.05,434.5,1,51,30,19.74,3263,1,San Mateo,0,0,Fiber Optic,37.556634,-122.317723,0,82.212,0,0,None,23393,0,1,0,0,6,3,130.0,118.44,0.0,434.5,0,0,94402
938,0,0,1,0,65,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),108.05,7118.9,0,32,15,41.34,6047,0,San Mateo,1,0,DSL,37.538309000000005,-122.305109,1,108.05,0,6,Offer B,37926,1,0,1,1,65,1,1068.0,2687.100000000001,0.0,7118.9,0,0,94403
939,0,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,320.45,0,46,0,2.74,3366,0,San Mateo,0,0,NA,37.556094,-122.27243700000001,0,19.9,0,0,None,31882,0,0,0,0,15,0,0.0,41.1,0.0,320.45,0,0,94404
940,0,0,0,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),21.05,531.55,0,55,0,47.31,2050,0,Alameda,0,0,NA,37.774633,-122.27443400000001,0,21.05,0,0,None,58555,0,0,0,0,24,3,0.0,1135.44,0.0,531.55,0,0,94501
941,0,0,0,1,13,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,30.15,382.2,0,50,19,0.0,3540,0,Alameda,0,0,DSL,37.724817,-122.22436299999998,0,30.15,2,0,None,13996,0,0,0,0,13,1,73.0,0.0,0.0,382.2,0,0,94502
942,1,0,0,0,24,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),79.85,2001,0,23,41,35.3,5128,0,Danville,0,1,DSL,37.791481,-121.903253,0,79.85,0,0,None,19777,0,0,0,1,24,0,0.0,847.1999999999998,0.0,2001.0,1,1,94506
943,0,0,1,0,72,0,No phone service,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),65.5,4919.7,0,56,4,0.0,4119,0,Alamo,1,0,Fiber Optic,37.855717,-121.994813,1,65.5,0,6,None,15187,1,1,1,1,72,1,0.0,0.0,0.0,4919.7,0,1,94507
944,0,0,1,1,54,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),104.1,5645.8,0,62,76,42.35,5795,0,Angwin,0,0,DSL,38.542448,-122.419923,1,104.1,3,3,Offer B,3641,0,0,1,1,54,2,4291.0,2286.9,0.0,5645.8,0,0,94508
945,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),74.4,215.8,1,32,26,23.82,2054,1,Antioch,0,0,Fiber Optic,37.980057,-121.801599,0,77.376,0,0,None,90891,0,0,0,0,3,5,56.0,71.46000000000002,0.0,215.8,0,0,94509
946,1,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.5,77.6,0,39,0,3.63,5053,0,Benicia,0,1,NA,38.113533000000004,-122.11926000000001,1,20.5,2,4,None,25578,0,0,1,0,4,2,0.0,14.52,0.0,77.6,0,0,94510
947,0,1,1,1,32,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,91.35,2896.55,0,66,30,5.73,2965,0,Bethel Island,1,0,Cable,38.050558,-121.646924,1,91.35,1,9,Offer C,2379,0,0,1,0,32,0,869.0,183.36,26.98,2896.55,0,0,94511
948,1,1,0,0,35,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.05,3395.8,1,71,21,20.83,2074,1,Birds Landing,1,1,Cable,38.140719,-121.838298,0,103.012,0,0,None,138,0,1,0,0,35,5,0.0,729.05,0.0,3395.8,0,1,94512
949,1,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.5,759.35,0,42,0,47.33,2009,0,Brentwood,0,1,NA,37.908242,-121.682472,1,20.5,1,8,None,26577,0,0,1,0,35,0,0.0,1656.55,0.0,759.35,0,0,94513
950,1,1,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.95,85.15,1,80,12,26.62,5900,1,Byron,0,1,Fiber Optic,37.83323,-121.60146100000001,0,46.74800000000001,0,0,Offer E,10153,0,2,0,0,2,5,10.0,53.24,0.0,85.15,0,0,94514
951,0,0,0,0,8,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,75.6,535.55,0,64,17,11.2,2934,0,Calistoga,0,0,DSL,38.629618,-122.593216,0,75.6,0,0,Offer E,7384,0,1,0,0,8,1,0.0,89.6,0.0,535.55,0,1,94515
952,1,0,0,0,22,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,55.1,1253.15,0,62,15,37.11,2729,0,Clayton,0,1,Fiber Optic,37.881842,-121.84811100000002,0,55.1,0,0,None,14239,1,0,0,0,22,1,0.0,816.42,0.0,1253.15,0,1,94517
953,0,0,0,0,15,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,58.95,955.15,0,57,11,30.54,4497,0,Concord,1,0,Cable,37.950247999999995,-122.02245500000001,0,58.95,0,0,None,27394,1,0,0,0,15,0,105.0,458.1,0.0,955.15,0,0,94518
954,1,0,0,0,22,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.1,2162.6,0,39,17,11.15,3729,0,Concord,0,1,Fiber Optic,37.990118,-122.012188,0,95.1,0,0,None,18650,0,0,0,1,22,2,0.0,245.3,0.0,2162.6,0,1,94519
955,1,0,1,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),44.7,44.7,1,21,80,32.08,3700,1,Concord,0,1,Fiber Optic,38.013825,-122.039144,1,46.48800000000001,0,1,None,36186,0,0,1,1,1,2,0.0,32.08,0.0,44.7,1,0,94520
956,0,0,1,1,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.45,1813.35,0,33,0,4.15,4993,0,Concord,0,0,NA,37.971421,-121.97150400000001,1,25.45,2,0,Offer A,39888,0,0,0,0,71,0,0.0,294.6500000000001,0.0,1813.35,0,0,94521
957,1,0,0,0,4,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,56.75,245.15,0,26,47,34.69,2401,0,Pleasant Hill,1,1,Fiber Optic,37.953379999999996,-122.07688600000002,0,56.75,0,0,Offer E,32685,0,0,0,0,4,2,0.0,138.76,0.0,245.15,1,1,94523
958,1,0,0,0,25,1,1,DSL,1,1,0,1,Month-to-month,0,Bank transfer (automatic),81.75,2028.8,0,59,23,25.2,5917,0,Crockett,1,1,DSL,38.049292,-122.22841499999998,0,81.75,0,0,None,3193,1,1,0,1,25,1,467.0,630.0,0.0,2028.8,0,0,94525
959,0,0,1,1,32,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,86.1,2723.75,0,45,57,26.66,4970,0,Danville,0,0,Cable,37.815459000000004,-121.977203,1,86.1,3,7,None,32873,0,0,1,0,32,1,0.0,853.12,0.0,2723.75,0,1,94526
960,1,1,1,0,7,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),29.8,220.45,0,80,13,0.0,2587,0,El Cerrito,0,1,DSL,37.924838,-122.28914499999999,1,29.8,0,10,Offer E,23141,0,0,1,0,7,0,2.87,0.0,11.83,220.45,0,1,94530
961,1,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.5,365.8,0,41,0,42.66,2259,0,Fairfield,0,1,NA,38.287136,-122.02711000000001,0,20.5,0,0,None,77683,0,0,0,0,17,2,0.0,725.2199999999998,0.0,365.8,0,0,94533
962,1,1,1,0,8,1,0,DSL,1,0,1,0,Month-to-month,0,Bank transfer (automatic),60.9,551.95,0,76,23,22.4,2136,0,Travis Afb,0,1,DSL,38.265899,-121.93946100000001,1,60.9,0,9,Offer E,9978,0,1,1,0,8,1,0.0,179.2,16.58,551.95,0,1,94535
963,0,1,0,0,56,1,1,DSL,1,0,0,1,Two year,0,Bank transfer (automatic),73.25,4054.2,0,80,8,37.3,4011,0,Fremont,1,0,DSL,37.572272999999996,-121.964583,0,73.25,0,0,None,66543,1,0,0,0,56,0,324.0,2088.8,17.16,4054.2,0,0,94536
964,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.7,45.7,1,36,19,10.41,3571,1,Fremont,0,1,Cable,37.505767999999996,-121.96247199999999,0,47.52800000000001,0,0,None,56126,0,0,0,0,1,4,0.0,10.41,0.0,45.7,0,0,94538
965,1,1,0,0,8,1,0,Fiber optic,1,0,1,1,Month-to-month,0,Credit card (automatic),100.3,832.35,1,66,30,11.57,5084,1,Fremont,0,1,DSL,37.516791,-121.89911699999999,0,104.31200000000001,0,0,None,46917,1,5,0,1,8,2,250.0,92.56,0.0,832.35,0,0,94539
966,1,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.25,112.3,1,53,0,9.14,4489,1,Hayward,0,1,NA,37.674002,-122.076796,0,19.25,0,0,None,60274,0,0,0,0,7,4,0.0,63.98,0.0,112.3,0,0,94541
967,1,0,0,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.85,60.65,0,50,0,19.58,5868,0,Hayward,0,1,NA,37.656695,-122.04836100000001,0,20.85,3,0,None,11147,0,2,0,0,3,1,0.0,58.74,0.0,60.65,0,0,94542
968,0,0,0,0,71,1,0,DSL,1,1,1,0,Two year,0,Credit card (automatic),77.35,5550.1,0,48,28,18.2,4846,0,Hayward,1,0,Fiber Optic,37.639215,-122.037554,0,77.35,0,0,Offer A,72993,1,0,0,0,71,0,0.0,1292.2,0.0,5550.1,0,1,94544
969,0,0,0,0,2,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.0,174.8,1,57,31,48.34,3391,1,Hayward,0,0,Fiber Optic,37.62984,-122.120843,0,99.84,0,0,None,27311,0,0,0,1,2,0,54.0,96.68,0.0,174.8,0,0,94545
970,0,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,90.55,90.55,1,30,56,15.44,2627,1,Castro Valley,0,0,DSL,37.708327000000004,-122.083473,0,94.17200000000001,0,0,Offer E,41698,0,0,0,1,1,5,0.0,15.44,0.0,90.55,0,0,94546
971,1,0,1,0,49,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Bank transfer (automatic),93.85,4733.1,0,30,26,47.17,5698,0,Hercules,0,1,Fiber Optic,37.991259,-122.214945,1,93.85,0,1,Offer B,22479,0,0,1,0,49,0,0.0,2311.33,0.0,4733.1,0,1,94547
972,1,0,0,0,58,1,0,DSL,0,1,1,0,Two year,0,Bank transfer (automatic),70.1,4048.95,0,26,69,47.47,4474,0,Lafayette,1,1,DSL,37.907777,-122.12716100000002,0,70.1,0,0,Offer B,23996,1,0,0,0,58,2,2794.0,2753.26,0.0,4048.95,1,0,94549
973,1,1,1,0,44,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,30.35,1359.7,1,73,31,0.0,4829,1,Livermore,0,1,Cable,37.571748,-121.65956200000001,1,31.564000000000004,0,2,None,75929,0,4,1,0,44,4,422.0,0.0,0.0,1359.7,0,0,94550
974,0,0,1,1,59,1,0,DSL,0,1,1,1,Two year,1,Credit card (automatic),75.95,4542.35,0,40,22,8.28,5446,0,Castro Valley,0,0,DSL,37.722727,-122.02157,1,75.95,0,4,Offer B,13212,1,0,1,1,59,1,999.0,488.52,0.0,4542.35,0,0,94552
975,1,0,0,0,71,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,108.05,7532.15,1,30,58,49.42,5200,1,Martinez,1,1,Cable,38.014457,-122.11543200000001,0,112.37200000000001,0,0,Offer A,46677,1,1,0,1,71,4,4369.0,3508.82,0.0,7532.15,0,0,94553
976,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.9,69.9,1,51,31,45.66,5367,1,Fremont,0,1,Cable,37.555473,-122.080312,0,72.69600000000001,0,0,Offer E,33883,0,0,0,0,1,2,0.0,45.66,0.0,69.9,0,0,94555
977,0,0,0,0,11,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.25,888.65,0,34,23,33.79,5902,0,Moraga,0,0,DSL,37.827946000000004,-122.10718500000002,0,75.25,0,0,Offer D,16510,0,0,0,0,11,2,0.0,371.69,0.0,888.65,0,1,94556
978,1,1,1,0,62,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,103.75,6383.35,1,77,18,7.11,5052,1,Napa,1,1,Fiber Optic,38.489789,-122.27011,1,107.9,0,1,None,63947,0,2,1,1,62,1,1149.0,440.82,0.0,6383.35,0,0,94558
979,0,0,1,1,35,1,0,DSL,1,0,0,0,One year,1,Bank transfer (automatic),54.95,1916,0,20,59,42.18,4858,0,Napa,0,0,Fiber Optic,38.232389000000005,-122.32494399999999,1,54.95,0,5,None,26894,1,0,1,0,35,0,1130.0,1476.3,0.0,1916.0,1,0,94559
980,0,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.5,413,0,23,0,10.97,5409,0,Newark,0,0,NA,37.504133,-122.032347,0,19.5,0,0,Offer D,42491,0,0,0,0,20,1,0.0,219.4,0.0,413.0,1,0,94560
981,1,0,1,1,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.6,808.95,0,21,0,22.96,2630,0,Oakley,0,1,NA,37.999406,-121.686241,1,19.6,1,9,Offer B,27607,0,0,1,0,40,0,0.0,918.4,0.0,808.95,1,0,94561
982,0,0,0,0,39,1,0,DSL,1,0,0,0,One year,1,Electronic check,47.85,1886.4,0,22,82,25.33,5531,0,Orinda,0,0,Cable,37.873915999999994,-122.20522,0,47.85,0,0,None,17964,0,0,0,0,39,1,1547.0,987.87,0.0,1886.4,1,0,94563
983,1,0,0,0,1,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.6,86.6,1,41,20,5.43,5228,1,Pinole,0,1,Fiber Optic,37.996462,-122.29371599999999,0,90.064,0,0,Offer E,16717,0,0,0,1,1,0,0.0,5.43,0.0,86.6,0,0,94564
984,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),23.75,1679.25,0,62,0,21.14,4923,0,Pittsburg,0,0,NA,38.006046999999995,-121.91683400000001,1,23.75,1,7,Offer A,78816,0,0,1,0,72,2,0.0,1522.08,0.0,1679.25,0,0,94565
985,0,1,1,0,33,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.6,2656.5,1,76,16,33.19,3601,1,Pleasanton,0,0,DSL,37.633361,-121.86239499999999,1,83.824,0,1,None,36669,0,0,1,0,33,2,0.0,1095.27,0.0,2656.5,0,1,94566
986,0,0,0,0,12,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),43.8,540.95,0,54,17,6.56,5706,0,Pope Valley,0,0,Fiber Optic,38.672708,-122.40321899999999,0,43.8,0,0,Offer D,494,0,0,0,0,12,0,0.0,78.72,0.0,540.95,0,1,94567
987,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.75,19.75,0,48,0,5.32,3595,0,Dublin,0,1,NA,37.713926,-121.928425,0,19.75,0,0,Offer E,29636,0,0,0,0,1,1,0.0,5.32,0.0,19.75,0,0,94568
988,1,0,0,1,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.15,537.35,0,20,0,30.36,4004,0,Port Costa,0,1,NA,38.035707,-122.196821,0,19.15,2,0,None,173,0,0,0,0,27,2,0.0,819.72,0.0,537.35,1,0,94569
989,1,0,1,1,34,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.6,678.8,0,53,0,26.03,4669,0,Rio Vista,0,1,NA,38.148862,-121.737696,1,19.6,0,7,None,5246,0,1,1,0,34,2,0.0,885.02,0.0,678.8,0,0,94571
990,0,0,1,0,56,1,0,Fiber optic,1,0,0,0,Two year,0,Bank transfer (automatic),80.3,4513.65,0,56,15,4.24,6203,0,Rodeo,1,0,DSL,38.027218,-122.23463000000001,1,80.3,0,9,Offer B,8506,0,0,1,0,56,0,677.0,237.44,0.0,4513.65,0,0,94572
991,0,0,0,0,58,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.35,1423.85,0,31,0,38.62,6190,0,Saint Helena,0,0,NA,38.581354,-122.296283,0,24.35,0,0,Offer B,9423,0,0,0,0,58,2,0.0,2239.96,0.0,1423.85,0,0,94574
992,0,0,1,1,22,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.25,555.4,0,30,0,25.98,4386,0,Deer Park,0,0,NA,38.554383,-122.474773,1,25.25,3,9,Offer D,223,0,0,1,0,22,1,0.0,571.5600000000002,0.0,555.4,0,0,94576
993,0,0,1,1,10,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),26.1,225.55,0,27,0,18.57,3179,0,San Leandro,0,0,NA,37.717196,-122.15933799999999,1,26.1,2,10,Offer D,41871,0,0,1,0,10,1,0.0,185.7,0.0,225.55,1,0,94577
994,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.0,268.45,0,23,0,1.61,3037,0,San Leandro,0,1,NA,37.704384000000005,-122.126703,0,20.0,0,0,Offer D,36568,0,0,0,0,13,2,0.0,20.93,0.0,268.45,1,0,94578
995,0,0,0,0,35,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Credit card (automatic),85.3,2917.5,1,28,45,45.14,2455,1,San Leandro,0,0,Cable,37.687264,-122.15728,0,88.712,0,0,Offer C,19815,1,2,0,1,35,6,1313.0,1579.9,23.89,2917.5,1,0,94579
996,0,0,0,0,34,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),70.0,2416.1,1,61,23,4.66,2318,1,San Lorenzo,0,0,Cable,37.676249,-122.132415,0,72.8,0,0,Offer C,26240,0,2,0,0,34,4,556.0,158.44,11.0,2416.1,0,0,94580
997,0,1,0,0,4,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.3,424.45,1,65,25,49.5,5419,1,San Ramon,0,0,Cable,37.766556,-121.97678400000001,0,98.072,0,0,Offer E,44078,0,0,0,1,4,0,106.0,198.0,0.0,424.45,0,0,94583
998,1,0,1,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.7,1492.1,0,19,0,21.72,6317,0,Suisun City,0,1,NA,38.197907,-122.01725800000001,1,20.7,0,1,Offer A,39279,0,0,1,0,72,1,0.0,1563.84,0.0,1492.1,1,0,94585
999,1,0,0,0,2,1,0,DSL,0,0,1,1,Month-to-month,0,Electronic check,70.3,132.4,0,21,48,23.52,4799,0,Sunol,0,1,DSL,37.587494,-121.86285600000001,0,70.3,0,0,None,790,1,0,0,1,2,1,64.0,47.04,0.0,132.4,1,0,94586
1000,0,0,0,0,7,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.35,660.9,1,46,16,48.36,3077,1,Union City,1,0,Cable,37.59485,-122.051521,0,99.164,0,0,Offer E,66472,0,0,0,1,7,1,106.0,338.52,34.29,660.9,0,0,94587
1001,1,1,1,0,27,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.5,1893.95,1,75,25,10.6,2377,1,Pleasanton,0,1,Cable,37.685052,-121.91206100000001,1,78.52,0,1,None,28568,0,3,1,0,27,1,473.0,286.2,0.0,1893.95,0,0,94588
1002,1,0,1,1,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.55,284.9,0,42,23,37.23,3708,0,Vallejo,0,1,DSL,38.161321,-122.271588,1,69.55,1,1,None,42209,0,0,1,0,4,1,66.0,148.92,0.0,284.9,0,0,94589
1003,0,0,0,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.85,784.25,0,28,0,26.49,3408,0,Vallejo,0,0,NA,38.104704999999996,-122.24738700000002,0,19.85,0,0,None,37218,0,0,0,0,37,1,0.0,980.13,0.0,784.25,1,0,94590
1004,1,0,0,0,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,417.7,0,59,0,34.39,2366,0,Vallejo,0,1,NA,38.105733,-122.18633799999999,0,20.0,0,0,Offer D,51665,0,0,0,0,21,0,0.0,722.19,0.0,417.7,0,0,94591
1005,0,1,1,0,53,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),95.85,5016.25,0,69,12,30.09,5325,0,Vallejo,0,0,Fiber Optic,38.093701,-122.27658899999999,1,95.85,0,1,None,159,0,0,1,0,53,1,0.0,1594.77,18.85,5016.25,0,1,94592
1006,0,0,0,0,18,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,90.1,1612.75,1,33,21,34.21,4260,1,Walnut Creek,0,0,Fiber Optic,37.862128000000006,-122.075197,0,93.704,0,0,None,18024,1,1,0,1,18,3,0.0,615.78,48.26,1612.75,0,1,94595
1007,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,68.95,119.75,1,26,43,30.73,5225,1,Walnut Creek,0,0,Cable,37.900662,-122.05278200000001,0,71.708,0,0,None,40917,0,2,0,1,2,2,51.0,61.46,0.0,119.75,1,0,94596
1008,1,0,1,1,32,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Credit card (automatic),99.55,3204.65,1,39,29,33.57,5026,1,Walnut Creek,0,1,Fiber Optic,37.916647999999995,-122.00848300000001,1,103.53200000000001,0,1,Offer C,26022,0,0,1,1,32,0,929.0,1074.24,35.82,3204.65,0,0,94598
1009,1,1,1,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,20.75,485.2,0,69,0,45.83,3418,0,Yountville,0,1,NA,38.421458,-122.365048,1,20.75,0,2,None,2873,0,0,1,0,23,1,0.0,1054.09,37.64,485.2,0,0,94599
1010,1,0,0,0,3,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,50.15,160.85,0,20,59,17.42,2085,0,Oakland,0,1,Cable,37.776523,-122.219268,0,50.15,0,0,None,54876,0,0,0,0,3,0,95.0,52.26000000000001,0.0,160.85,1,0,94601
1011,0,0,1,1,71,0,No phone service,DSL,1,1,1,1,Two year,0,Mailed check,58.65,4145.25,0,31,8,0.0,4151,0,Oakland,0,0,Fiber Optic,37.803883,-122.208417,1,58.65,0,3,Offer A,28900,1,0,1,1,71,1,332.0,0.0,0.0,4145.25,0,0,94602
1012,1,0,0,0,9,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.9,827.45,0,41,3,30.8,5017,0,Oakland,0,1,DSL,37.739113,-122.175602,0,95.9,0,0,None,31392,1,0,0,1,9,0,25.0,277.2,0.0,827.45,0,0,94603
1013,0,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,49.5,49.5,0,56,8,16.99,5262,0,Oakland,0,0,Fiber Optic,37.758019,-122.138678,0,49.5,0,0,None,42854,0,1,0,0,1,2,0.0,16.99,0.0,49.5,0,0,94605
1014,1,0,1,1,18,1,0,DSL,0,0,0,1,Month-to-month,0,Electronic check,57.45,990.85,1,53,24,2.86,2989,1,Oakland,1,1,DSL,37.792489,-122.24431399999999,1,59.74800000000001,0,1,None,41876,0,1,1,1,18,4,0.0,51.48,15.73,990.85,0,1,94606
1015,1,0,1,1,12,1,0,DSL,0,0,0,1,One year,0,Credit card (automatic),53.65,696.35,1,27,29,27.82,2595,1,Oakland,0,1,Fiber Optic,37.80707,-122.29740100000001,1,55.79600000000001,0,1,None,21054,0,1,1,1,12,2,0.0,333.8400000000001,0.0,696.35,1,1,94607
1016,1,0,1,0,71,1,1,DSL,1,1,0,1,Two year,1,Mailed check,80.1,5585.4,0,36,20,10.97,6045,0,Emeryville,1,1,Fiber Optic,37.83726,-122.287648,1,80.1,0,5,Offer A,24589,1,0,1,1,71,1,111.71,778.87,0.0,5585.4,0,1,94608
1017,0,0,0,0,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),24.4,1601.2,0,36,0,15.93,5887,0,Oakland,0,0,NA,37.834340999999995,-122.26437,0,24.4,0,0,Offer B,21097,0,0,0,0,64,1,0.0,1019.52,0.0,1601.2,0,0,94609
1018,1,0,0,0,4,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,40.05,162.45,0,33,13,0.0,2664,0,Oakland,0,1,Fiber Optic,37.808731,-122.238708,0,40.05,0,0,None,29964,1,0,0,1,4,0,21.0,0.0,0.0,162.45,0,0,94610
1019,0,0,0,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.5,470.2,0,33,0,13.98,5652,0,Oakland,0,0,NA,37.828416,-122.21600500000001,0,19.5,0,0,Offer D,36517,0,0,0,0,23,3,0.0,321.54,0.0,470.2,0,0,94611
1020,0,0,1,1,39,1,0,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),51.05,2066,0,59,11,15.06,3154,0,Oakland,0,0,DSL,37.809014000000005,-122.26973899999999,1,51.05,2,3,None,11702,0,0,1,0,39,1,227.0,587.34,0.0,2066.0,0,0,94612
1021,1,0,1,0,28,1,0,DSL,1,0,0,0,One year,0,Mailed check,54.35,1426.45,0,27,48,33.63,5105,0,Oakland,0,1,Cable,37.84551,-122.23518100000001,1,54.35,0,1,None,15438,1,0,1,0,28,1,0.0,941.64,0.0,1426.45,1,1,94618
1022,0,1,0,0,5,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,84.7,392.5,0,73,4,14.22,2660,0,Oakland,0,0,Fiber Optic,37.787186,-122.14633,0,84.7,0,0,Offer E,24518,0,1,0,0,5,1,0.0,71.10000000000002,41.2,392.5,0,1,94619
1023,0,1,1,0,45,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.1,3861.45,0,67,24,40.85,2701,0,Oakland,1,0,Cable,37.750553000000004,-122.197175,1,86.1,0,5,None,30751,0,0,1,0,45,0,0.0,1838.25,12.19,3861.45,0,1,94621
1024,1,0,0,0,37,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.35,2552.9,0,62,25,28.84,5402,0,Berkeley,0,1,DSL,37.866009000000005,-122.28622800000001,0,70.35,0,0,None,15638,0,0,0,0,37,1,0.0,1067.08,0.0,2552.9,0,1,94702
1025,0,1,1,0,60,1,0,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),110.0,6668.35,0,69,30,24.62,4953,0,Berkeley,1,0,Fiber Optic,37.863843,-122.27568400000001,1,110.0,0,2,None,19763,1,0,1,0,60,1,0.0,1477.2,0.0,6668.35,0,1,94703
1026,1,1,0,0,8,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.6,819.4,1,75,32,40.45,5906,1,Berkeley,1,1,Cable,37.871415999999996,-122.246597,0,104.624,0,0,Offer E,21205,0,0,0,0,8,4,0.0,323.6,0.0,819.4,0,1,94704
1027,0,0,0,0,47,1,1,Fiber optic,1,0,1,0,One year,0,Credit card (automatic),94.9,4615.25,0,30,69,40.25,4510,0,Berkeley,1,0,DSL,37.858897999999996,-122.24051200000001,0,94.9,0,0,Offer B,12448,0,0,0,0,47,0,3185.0,1891.75,0.0,4615.25,0,0,94705
1028,1,0,1,1,26,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,83.75,2070.6,1,62,29,35.9,2404,1,Albany,0,1,DSL,37.890274,-122.29519199999999,1,87.10000000000002,0,1,Offer C,15882,0,1,1,0,26,1,600.0,933.4,0.0,2070.6,0,0,94706
1029,0,1,1,1,3,1,0,Fiber optic,1,0,1,0,Month-to-month,1,Mailed check,88.3,273.75,1,68,2,25.77,4486,1,Berkeley,0,0,DSL,37.897753,-122.27939099999999,1,91.83200000000001,0,1,Offer E,11889,1,0,1,0,3,2,5.0,77.31,0.0,273.75,0,0,94707
1030,0,0,1,1,50,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.75,3557.7,0,39,23,10.21,4539,0,Berkeley,0,0,Fiber Optic,37.897743,-122.263124,1,69.75,3,8,Offer B,10737,0,0,1,0,50,0,818.0,510.50000000000006,0.0,3557.7,0,0,94708
1031,1,0,1,1,27,1,1,DSL,0,0,1,1,Month-to-month,0,Bank transfer (automatic),71.6,1957.1,0,30,59,13.55,3773,0,Berkeley,0,1,Fiber Optic,37.878554,-122.26608999999999,1,71.6,2,1,None,10147,1,0,1,1,27,1,0.0,365.85,0.0,1957.1,0,1,94709
1032,0,1,0,0,8,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,92.1,729.95,1,71,10,42.93,5662,1,Berkeley,1,0,Cable,37.872902,-122.30370800000001,0,95.784,0,0,Offer E,8157,0,0,0,0,8,0,0.0,343.44,0.0,729.95,0,1,94710
1033,0,0,1,0,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),23.65,1416.75,0,49,0,8.91,4671,0,Richmond,0,0,NA,37.945288,-122.383941,1,23.65,0,4,None,28450,0,2,1,0,62,1,0.0,552.42,0.0,1416.75,0,0,94801
1034,0,0,1,0,71,1,0,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),81.85,5924.4,0,25,58,6.23,4090,0,El Sobrante,1,0,Fiber Optic,37.963995000000004,-122.288296,1,81.85,0,4,Offer A,25399,1,0,1,1,71,0,0.0,442.33,0.0,5924.4,1,1,94803
1035,1,0,0,0,66,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.1,1697.7,0,39,0,49.13,6025,0,Richmond,0,1,NA,37.921034000000006,-122.341798,0,25.1,0,0,Offer A,39089,0,0,0,0,66,0,0.0,3242.580000000001,0.0,1697.7,0,0,94804
1036,1,0,1,1,68,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.7,7849.85,0,61,24,32.59,5671,0,Richmond,1,1,Fiber Optic,37.941456,-122.320968,1,114.7,1,5,Offer A,13984,1,0,1,1,68,0,0.0,2216.120000000001,0.0,7849.85,0,1,94805
1037,0,0,0,0,13,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Electronic check,49.15,649.4,0,47,27,0.0,3000,0,San Pablo,1,0,DSL,37.980269,-122.34263500000002,0,49.15,0,0,Offer D,55720,0,0,0,1,13,1,0.0,0.0,0.0,649.4,0,1,94806
1038,1,0,1,0,56,1,0,Fiber optic,0,0,0,1,One year,1,Electronic check,80.9,4557.5,0,37,24,46.18,5344,0,San Rafael,0,1,Cable,37.972662,-122.491452,1,80.9,0,3,None,40239,0,0,1,1,56,1,0.0,2586.08,0.0,4557.5,0,1,94901
1039,1,0,1,0,38,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,79.45,3013.05,1,44,14,35.61,2405,1,San Rafael,0,1,Cable,38.018065,-122.546024,1,82.62799999999999,0,1,None,28403,0,1,1,0,38,4,422.0,1353.18,9.36,3013.05,0,0,94903
1040,1,1,0,0,14,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Credit card (automatic),90.45,1266.1,1,74,26,11.31,4777,1,Greenbrae,0,1,DSL,37.946616999999996,-122.563571,0,94.068,0,0,None,12010,0,0,0,0,14,0,329.0,158.34,0.0,1266.1,0,0,94904
1041,0,0,0,1,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.3,360.35,0,56,0,44.05,2870,0,Belvedere Tiburon,0,0,NA,37.885628999999994,-122.46858,0,19.3,0,0,Offer D,13065,0,0,0,0,16,1,0.0,704.8,0.0,360.35,0,0,94920
1042,0,0,1,1,14,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.2,1046.5,0,60,17,23.0,5819,0,Bodega,0,0,Cable,38.343282,-122.9755,1,70.2,2,0,Offer D,584,0,0,0,0,14,0,0.0,322.0,0.0,1046.5,0,1,94922
1043,1,0,1,1,32,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.75,2347.9,1,37,6,5.99,2356,1,Bodega Bay,0,1,Cable,38.377165000000005,-123.037957,1,72.54,0,1,None,1785,0,0,1,0,32,3,0.0,191.68,19.67,2347.9,0,1,94923
1044,0,0,0,0,8,1,0,DSL,1,0,0,0,One year,0,Bank transfer (automatic),54.25,447.75,0,37,27,42.78,2237,0,Bolinas,0,0,DSL,37.943087,-122.72379,0,54.25,0,0,None,1573,1,0,0,0,8,0,0.0,342.24,0.0,447.75,0,1,94924
1045,0,0,1,1,43,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),99.3,4209.95,0,29,59,5.25,3280,0,Corte Madera,1,0,Fiber Optic,37.924014,-122.51169399999999,1,99.3,2,8,None,9038,0,2,1,1,43,3,0.0,225.75,0.0,4209.95,1,1,94925
1046,0,0,0,0,52,1,1,DSL,1,0,1,0,One year,0,Credit card (automatic),74.0,3877.65,0,31,21,21.38,5806,0,Rohnert Park,1,0,Fiber Optic,38.347190000000005,-122.697822,0,74.0,0,0,None,42544,1,0,0,0,52,0,81.43,1111.76,0.0,3877.65,0,1,94928
1047,1,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.25,152.3,0,35,21,28.19,2166,0,Dillon Beach,0,1,Fiber Optic,38.24458,-122.956268,0,50.25,0,0,None,330,1,0,0,0,3,0,0.0,84.57000000000002,0.0,152.3,0,1,94929
1048,1,0,0,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.8,572.2,0,42,0,46.12,5696,0,Fairfax,0,1,NA,37.971751,-122.611873,0,19.8,0,0,None,8486,0,0,0,0,29,3,0.0,1337.48,0.0,572.2,0,0,94930
1049,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,19.65,1,50,0,6.08,5881,1,Cotati,0,0,NA,38.326215000000005,-122.71874199999999,0,19.65,0,0,Offer E,7936,0,0,0,0,1,0,0.0,6.08,0.0,19.65,0,0,94931
1050,1,1,0,0,12,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,43.65,526.95,1,77,11,0.0,2437,1,Forest Knolls,1,1,Cable,38.010092,-122.68944199999999,0,45.396,0,0,None,1025,1,4,0,0,12,2,58.0,0.0,0.0,526.95,0,0,94933
1051,0,0,1,1,16,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Credit card (automatic),35.5,552.7,0,48,53,0.0,2069,0,Inverness,0,0,Cable,38.099323,-122.945723,1,35.5,3,1,Offer D,1004,0,0,1,1,16,2,0.0,0.0,0.0,552.7,0,1,94937
1052,0,0,0,0,40,1,1,DSL,0,0,1,1,One year,1,Mailed check,80.75,3208.65,0,41,19,33.83,2047,0,Lagunitas,1,0,Fiber Optic,38.021772,-122.691744,0,80.75,0,0,None,821,1,0,0,1,40,1,610.0,1353.1999999999996,0.0,3208.65,0,0,94938
1053,0,0,0,0,5,0,No phone service,DSL,0,0,0,1,Month-to-month,0,Electronic check,39.5,210.75,1,55,2,0.0,2863,1,Larkspur,1,0,Cable,37.937082000000004,-122.53236899999999,0,41.08,0,0,Offer E,6773,0,0,0,1,5,4,4.0,0.0,39.27,210.75,0,0,94939
1054,1,0,1,0,40,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),97.1,3706.95,1,58,25,16.33,3099,1,Marshall,0,1,DSL,38.129308,-122.83481499999999,1,100.984,0,1,Offer B,406,0,0,1,1,40,2,927.0,653.1999999999998,41.85,3706.95,0,0,94940
1055,0,0,0,0,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.55,620.75,0,47,0,41.33,2691,0,Mill Valley,0,0,NA,37.901371000000005,-122.572024,0,19.55,0,0,None,28727,0,0,0,0,36,0,0.0,1487.88,0.0,620.75,0,0,94941
1056,0,0,0,0,5,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.0,412.5,1,26,46,43.99,3937,1,Novato,0,0,DSL,38.135897,-122.56368300000001,0,83.2,0,0,Offer E,16429,0,0,0,1,5,0,0.0,219.95,40.0,412.5,1,1,94945
1057,0,0,0,0,10,1,0,Fiber optic,1,0,1,0,Month-to-month,1,Mailed check,84.7,832.05,1,40,20,45.69,5686,1,Nicasio,0,0,Cable,38.065359,-122.665566,0,88.08800000000002,0,0,None,607,0,0,0,0,10,0,166.0,456.9,12.81,832.05,0,0,94946
1058,1,0,1,1,2,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),89.55,185.55,1,49,25,8.86,3851,1,Novato,0,1,Fiber Optic,38.112165999999995,-122.63438400000001,1,93.132,0,1,Offer E,24741,0,1,1,1,2,1,46.0,17.72,0.0,185.55,0,0,94947
1059,1,0,0,0,23,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,90.6,1943.2,1,21,76,38.69,4359,1,Novato,0,1,Cable,38.067204,-122.524004,0,94.22399999999999,0,0,None,13361,1,0,0,1,23,3,1477.0,889.8699999999999,4.73,1943.2,1,0,94949
1060,1,0,1,1,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.05,505.9,0,49,0,45.28,2403,0,Olema,0,1,NA,38.052209000000005,-122.775567,1,20.05,0,10,None,248,0,0,1,0,26,0,0.0,1177.28,0.0,505.9,0,0,94950
1061,0,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,112.4,8046.85,0,80,2,15.23,6144,0,Penngrove,1,0,Fiber Optic,38.325599,-122.642352,1,112.4,0,5,Offer A,3777,0,0,1,0,72,0,0.0,1096.56,0.0,8046.85,0,1,94951
1062,0,0,1,0,34,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),50.2,1815.3,0,33,7,40.67,4352,0,Petaluma,0,0,Cable,38.237018,-122.77871999999999,1,50.2,0,6,None,31930,1,0,1,0,34,1,127.0,1382.78,0.0,1815.3,0,0,94952
1063,1,0,0,0,10,1,0,DSL,1,0,1,0,Month-to-month,0,Bank transfer (automatic),62.25,612.95,0,32,17,7.65,3415,0,Petaluma,0,1,Fiber Optic,38.235021,-122.557332,0,62.25,0,0,Offer D,35419,1,1,0,0,10,1,104.0,76.5,0.0,612.95,0,0,94954
1064,0,0,0,0,14,1,0,DSL,1,0,0,0,One year,0,Mailed check,55.7,795.15,0,52,26,27.68,4978,0,Point Reyes Station,0,0,DSL,38.060264000000004,-122.830646,0,55.7,0,0,None,1885,1,0,0,0,14,1,207.0,387.52,0.0,795.15,0,0,94956
1065,0,0,0,0,23,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Bank transfer (automatic),90.05,2169.8,1,64,4,3.55,4650,1,San Anselmo,0,0,Fiber Optic,37.99272,-122.575026,0,93.652,0,0,None,16849,0,0,0,0,23,2,87.0,81.64999999999998,27.38,2169.8,0,0,94960
1066,1,0,1,0,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.65,973.1,0,63,0,6.54,2021,0,San Geronimo,0,1,NA,38.004740000000005,-122.66371699999999,1,19.65,0,7,None,548,0,0,1,0,47,1,0.0,307.38,0.0,973.1,0,0,94963
1067,1,0,1,0,24,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,89.25,2210.2,0,36,8,10.23,5436,0,San Quentin,0,1,Cable,37.942551,-122.491642,1,89.25,0,2,None,6448,1,0,1,1,24,0,0.0,245.52,0.0,2210.2,0,1,94964
1068,1,0,1,0,49,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),99.05,4853.75,1,54,24,20.48,5157,1,Sausalito,0,1,Fiber Optic,37.848641,-122.51569199999999,1,103.012,0,1,Offer B,11213,0,0,1,1,49,0,1165.0,1003.52,14.24,4853.75,0,0,94965
1069,1,1,0,0,20,1,0,DSL,1,0,0,0,One year,0,Mailed check,54.0,1055.9,0,68,21,22.31,5090,0,Stinson Beach,0,1,Fiber Optic,37.921137,-122.65756200000001,0,54.0,0,0,None,781,1,0,0,0,20,1,0.0,446.2,0.0,1055.9,0,1,94970
1070,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),69.75,144.55,1,46,26,26.44,5667,1,Tomales,0,0,Cable,38.240769,-122.90104099999999,0,72.54,0,0,None,384,0,4,0,0,2,2,3.76,52.88,0.0,144.55,0,1,94971
1071,0,0,0,0,2,1,0,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),49.05,91.1,1,42,14,14.7,2960,1,Valley Ford,0,0,Fiber Optic,38.339996,-122.935056,0,51.012,0,0,Offer E,66,0,2,0,0,2,1,13.0,29.4,0.0,91.1,0,0,94972
1072,1,0,0,0,22,0,No phone service,DSL,0,0,1,1,Two year,0,Bank transfer (automatic),56.75,1304.85,0,62,19,0.0,4574,0,Woodacre,1,1,DSL,38.005839,-122.638155,0,56.75,0,0,None,1449,1,0,0,1,22,1,0.0,0.0,0.0,1304.85,0,1,94973
1073,1,0,0,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),98.05,713,1,32,32,9.25,2561,1,Alviso,1,1,Cable,37.449537,-121.994813,0,101.97200000000001,0,0,Offer E,2147,0,1,0,1,7,3,228.0,64.75,0.0,713.0,0,0,95002
1074,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,21.1,21.1,0,31,0,18.81,2810,0,Aptos,0,1,NA,37.013471,-121.877877,0,21.1,0,0,None,24227,0,1,0,0,1,1,0.0,18.81,0.0,21.1,0,0,95003
1075,0,0,1,1,59,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),96.65,5580.8,0,35,53,48.07,5266,0,Aromas,0,0,Fiber Optic,36.878364000000005,-121.62978100000001,1,96.65,5,2,None,3373,1,0,1,1,59,0,2958.0,2836.13,0.0,5580.8,0,0,95004
1076,0,0,1,1,58,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),24.5,1497.9,0,44,0,36.45,4455,0,Ben Lomond,0,0,NA,37.078873,-122.09038600000001,1,24.5,0,9,None,6407,0,0,1,0,58,1,0.0,2114.100000000001,9.22,1497.9,0,0,95005
1077,0,0,0,0,41,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),114.5,4527.45,1,23,65,21.56,3038,1,Boulder Creek,1,0,DSL,37.171727000000004,-122.14296100000001,0,119.08,0,0,Offer B,10520,1,0,0,1,41,4,2943.0,883.9599999999998,0.0,4527.45,1,0,95006
1078,0,1,0,0,59,1,1,Fiber optic,0,1,0,0,Two year,1,Credit card (automatic),79.2,4590.35,0,71,2,6.13,5400,0,Brookdale,0,0,DSL,37.106902000000005,-122.10000600000001,0,79.2,0,0,None,1007,0,0,0,0,59,0,0.0,361.67,0.0,4590.35,0,1,95007
1079,0,0,1,1,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.55,200.2,0,61,19,1.67,5998,0,Campbell,0,0,Cable,37.279689000000005,-121.954567,1,69.55,2,3,None,44976,0,0,1,0,3,1,38.0,5.01,33.8,200.2,0,0,95008
1080,1,0,0,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.05,614.45,0,50,0,14.91,3398,0,Capitola,0,1,NA,36.977025,-121.95286399999999,0,20.05,0,0,None,9673,0,0,0,0,32,1,0.0,477.12,9.73,614.45,0,0,95010
1081,1,1,1,0,46,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.85,4564.9,0,74,22,4.2,2641,0,Castroville,1,1,Fiber Optic,36.784481,-121.759054,1,98.85,0,6,None,8582,0,0,1,0,46,1,100.43,193.2,0.0,4564.9,0,1,95012
1082,1,0,1,1,0,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.75, ,0,39,0,22.83,4950,0,Cupertino,0,1,NA,37.306612,-122.080621,1,25.75,1,5,None,54431,0,0,1,0,10,1,0.0,228.3,0.0,257.5,0,0,95014
1083,1,0,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.95,171.15,1,51,15,17.33,3533,1,Davenport,0,1,Fiber Optic,37.114335,-122.23716200000001,0,84.18799999999999,0,0,Offer E,857,0,0,0,1,2,0,26.0,34.66,0.0,171.15,0,0,95017
1084,0,0,1,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.6,1012.4,0,41,0,8.25,4848,0,Felton,0,0,NA,37.089110999999995,-122.06221299999999,1,19.6,0,0,None,8728,0,0,0,0,52,0,0.0,429.0,46.07,1012.4,0,0,95018
1085,0,1,0,0,13,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.3,940.35,1,73,23,40.37,2995,1,Freedom,1,0,DSL,36.936228,-121.785559,0,77.27199999999999,0,0,None,4753,0,2,0,0,13,1,216.0,524.81,0.0,940.35,0,0,95019
1086,0,1,0,0,11,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),89.7,1047.7,1,68,30,3.96,2202,1,Gilroy,0,0,Cable,37.03889,-121.52895500000001,0,93.288,0,0,None,49968,0,0,0,0,11,4,314.0,43.56,0.0,1047.7,0,0,95020
1087,1,0,0,0,32,1,1,Fiber optic,1,0,0,0,Month-to-month,0,Bank transfer (automatic),87.65,2766.4,0,53,25,6.2,2426,0,Escondido,0,1,DSL,33.141265000000004,-116.967221,0,87.65,0,0,None,48690,1,0,0,0,32,0,69.16,198.4,47.87,2766.4,0,1,92027
1088,1,1,1,0,17,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),100.45,1622.45,1,74,18,28.18,5508,1,Los Gatos,1,1,Cable,37.222842,-121.988727,1,104.46799999999999,0,1,None,13290,0,0,1,0,17,0,0.0,479.06,0.0,1622.45,0,1,95030
1089,0,0,0,0,16,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.75,1129.35,0,35,16,13.04,3574,0,Los Gatos,0,0,DSL,37.233034,-121.947427,0,74.75,0,0,None,24443,0,0,0,0,16,0,181.0,208.64,39.99,1129.35,0,0,95032
1090,0,0,0,0,51,1,1,Fiber optic,1,1,1,1,One year,0,Bank transfer (automatic),107.45,5680.9,0,62,6,7.54,5446,0,Los Gatos,1,0,Fiber Optic,37.160194,-121.94561100000001,0,107.45,0,0,None,10172,0,0,0,1,51,1,341.0,384.54,14.76,5680.9,0,0,95033
1091,1,0,0,0,29,1,0,DSL,0,0,1,1,One year,1,Bank transfer (automatic),75.35,2243.9,0,30,27,3.69,4422,0,Milpitas,1,1,Fiber Optic,37.441931,-121.878502,0,75.35,0,0,None,62848,1,0,0,1,29,1,60.59,107.01,2.24,2243.9,0,1,95035
1092,1,0,1,0,70,1,0,DSL,1,1,0,0,Two year,0,Credit card (automatic),64.95,4523.25,0,24,41,1.63,5669,0,Morgan Hill,1,1,Fiber Optic,37.161544,-121.649371,1,64.95,0,1,Offer A,41707,1,0,1,0,70,1,0.0,114.1,42.89,4523.25,1,1,95037
1093,0,0,1,1,71,1,1,Fiber optic,1,0,0,1,Two year,0,Electronic check,100.45,7159.7,0,25,59,32.16,6171,0,Moss Landing,1,0,Fiber Optic,36.863303,-121.781632,1,100.45,2,4,Offer A,899,1,0,1,1,71,0,422.42,2283.36,16.12,7159.7,1,1,95039
1094,1,0,1,1,41,1,1,DSL,0,1,1,0,One year,0,Bank transfer (automatic),68.5,2839.95,0,28,51,13.58,3877,0,Mount Hermon,1,1,Fiber Optic,37.051165999999995,-122.05619399999999,1,68.5,0,4,None,77,0,0,1,0,41,0,1448.0,556.78,38.37,2839.95,1,0,95041
1095,1,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.55,80.55,0,49,19,5.93,3154,0,Paicines,0,1,Fiber Optic,36.525703,-120.952122,0,80.55,0,0,None,813,0,0,0,0,1,0,0.0,5.93,0.0,80.55,0,0,95043
1096,0,0,1,0,7,1,0,DSL,1,0,1,1,Month-to-month,0,Bank transfer (automatic),81.25,580.1,0,38,9,12.16,5928,0,San Juan Bautista,1,0,DSL,36.810567999999996,-121.503022,1,81.25,0,4,None,3402,1,1,1,1,7,2,0.0,85.12,47.36,580.1,0,1,95045
1097,1,0,1,1,25,1,0,Fiber optic,0,0,1,1,One year,1,Electronic check,90.4,2178.6,1,63,4,35.27,5801,1,San Martin,0,1,Fiber Optic,37.084697,-121.606417,1,94.016,0,1,None,5671,0,0,1,1,25,0,87.0,881.7500000000001,0.0,2178.6,0,0,95046
1098,1,0,1,1,67,1,1,Fiber optic,1,1,0,0,One year,0,Electronic check,89.55,6038.55,0,60,11,18.29,6194,0,Santa Clara,0,1,DSL,37.351214,-121.952417,1,89.55,1,10,Offer A,36349,1,0,1,0,67,2,664.0,1225.4299999999996,33.76,6038.55,0,0,95050
1099,1,0,1,1,5,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,55.7,259.4,0,38,12,18.97,3598,0,Santa Clara,0,1,DSL,37.348129,-121.98468999999999,1,55.7,1,3,None,52986,1,0,1,0,5,0,31.0,94.85,0.0,259.4,0,0,95051
1100,1,0,0,1,15,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,24.8,324.15,0,53,0,32.54,3965,0,Santa Clara,0,1,NA,37.393553999999995,-121.96511399999999,0,24.8,3,0,None,13031,0,0,0,0,15,0,0.0,488.1,12.8,324.15,0,0,95054
1101,0,0,1,1,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.0,417.65,0,21,0,38.6,3402,0,Santa Cruz,0,0,NA,36.993451,-122.098858,1,20.0,3,4,None,43192,0,0,1,0,20,1,0.0,772.0,9.73,417.65,1,0,95060
1102,1,0,1,1,3,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,56.15,168.15,1,21,57,29.29,2539,1,Santa Cruz,1,1,Fiber Optic,36.974575,-121.991149,1,58.396,0,1,Offer E,36631,0,2,1,1,3,1,96.0,87.87,0.0,168.15,1,0,95062
1103,1,0,1,1,54,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,105.2,5637.85,0,50,57,7.25,5546,0,Santa Cruz,0,1,Cable,37.007882,-122.065975,1,105.2,3,9,None,4563,1,0,1,1,54,0,0.0,391.5,23.01,5637.85,0,1,95064
1104,1,0,0,0,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.55,839.4,0,32,0,48.41,5293,0,Santa Cruz,0,1,NA,37.031403999999995,-121.98186499999998,0,19.55,0,0,None,8365,0,0,0,0,42,0,0.0,2033.22,12.16,839.4,0,0,95065
1105,0,0,1,0,9,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.75,769.1,0,24,59,6.78,4654,0,Scotts Valley,0,0,Fiber Optic,37.070177,-122.010077,1,79.75,0,3,None,14574,0,0,1,1,9,0,0.0,61.02,0.0,769.1,1,1,95066
1106,0,0,0,0,63,1,1,Fiber optic,0,1,1,1,Two year,0,Bank transfer (automatic),97.45,6253,0,24,48,37.76,4769,0,Saratoga,0,0,Fiber Optic,37.257771999999996,-122.051824,0,97.45,0,0,None,30589,0,0,0,1,63,0,0.0,2378.88,0.0,6253.0,1,1,95070
1107,0,0,1,0,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.25,1641.8,0,57,0,39.78,4884,0,Soquel,0,0,NA,37.023669,-121.94646100000001,1,24.25,0,10,Offer A,9823,0,0,1,0,69,0,0.0,2744.82,45.75,1641.8,0,0,95073
1108,0,0,0,0,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.6,1678.05,0,24,0,36.5,5294,0,Watsonville,0,0,NA,36.931653999999995,-121.75238300000001,0,24.6,0,0,Offer A,81141,0,0,0,0,69,2,0.0,2518.5,28.42,1678.05,1,0,95076
1109,1,0,1,0,40,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,50.15,2058.5,0,32,28,24.3,2454,0,San Jose,0,1,Cable,37.34667,-121.91001899999999,1,50.15,0,7,None,18197,0,0,1,0,40,2,0.0,972.0,37.03,2058.5,0,1,95110
1110,1,0,0,0,60,0,No phone service,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),39.6,2424.5,0,38,25,0.0,5544,0,San Jose,1,1,DSL,37.284265000000005,-121.827673,0,39.6,0,0,Offer B,57748,0,0,0,0,60,0,60.61,0.0,38.46,2424.5,0,1,95111
1111,0,0,0,0,4,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Bank transfer (automatic),94.4,387.2,1,59,20,39.68,4249,1,San Jose,1,0,Fiber Optic,37.343827000000005,-121.883119,0,98.17600000000002,0,0,Offer E,52334,1,0,0,1,4,0,77.0,158.72,0.0,387.2,0,0,95112
1112,0,1,0,0,71,1,1,DSL,1,1,1,1,Two year,0,Mailed check,89.85,6293.45,0,69,22,37.39,4994,0,San Jose,1,0,Fiber Optic,37.333851,-121.891147,0,89.85,0,0,Offer A,561,1,0,0,0,71,2,0.0,2654.69,0.0,6293.45,0,1,95113
1113,0,0,1,0,37,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),78.95,2839.65,1,62,32,37.49,3982,1,San Jose,1,0,Cable,37.350284,-121.852855,1,82.10799999999999,0,0,None,51706,0,0,0,0,37,2,0.0,1387.13,0.0,2839.65,0,1,95116
1114,1,0,1,0,32,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),98.85,3145.9,0,33,9,47.89,3981,0,San Jose,0,1,Fiber Optic,37.311088,-121.961786,1,98.85,0,3,None,29914,0,0,1,1,32,0,28.31,1532.48,0.0,3145.9,0,1,95117
1115,1,0,0,0,39,1,1,DSL,0,0,0,0,Two year,1,Credit card (automatic),53.85,2200.7,0,60,16,5.4,2380,0,San Jose,0,1,Fiber Optic,37.255479,-121.88983799999998,0,53.85,0,0,None,31926,1,0,0,0,39,3,352.0,210.6,46.66,2200.7,0,0,95118
1116,0,0,0,0,38,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,24.25,914.4,0,36,0,46.18,2997,0,San Jose,0,0,NA,37.233226,-121.78809,0,24.25,0,0,None,10155,0,0,0,0,38,0,0.0,1754.84,35.61,914.4,0,0,95119
1117,1,0,0,0,52,1,1,Fiber optic,0,0,0,1,Two year,1,Credit card (automatic),89.45,4577.75,0,32,17,15.1,5386,0,San Jose,1,1,Fiber Optic,37.186141,-121.843554,0,89.45,0,0,Offer B,37090,0,0,0,1,52,0,778.0,785.1999999999998,18.89,4577.75,0,0,95120
1118,0,0,1,1,48,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),105.25,4997.5,0,57,53,30.41,4275,0,San Jose,0,0,Fiber Optic,37.304681,-121.809955,1,105.25,3,1,Offer B,37127,0,0,1,1,48,2,0.0,1459.68,1.66,4997.5,0,1,95121
1119,1,0,1,1,70,0,No phone service,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),59.5,4144.8,0,21,30,0.0,4031,0,San Jose,1,1,Fiber Optic,37.32886,-121.83456699999999,1,59.5,0,7,Offer A,59841,1,0,1,1,70,0,1243.0,0.0,23.72,4144.8,1,0,95122
1120,1,0,0,0,20,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),70.55,1493.55,0,56,26,3.8,5790,0,San Jose,0,1,Fiber Optic,37.238758000000004,-121.828375,0,70.55,0,0,None,59632,0,0,0,0,20,3,0.0,76.0,17.6,1493.55,0,1,95123
1121,0,0,0,0,50,1,1,DSL,1,0,1,1,One year,1,Credit card (automatic),82.5,4179.1,0,59,2,21.25,5258,0,San Jose,1,0,DSL,37.257063,-121.92303700000001,0,82.5,0,0,Offer B,45257,1,0,0,1,50,2,84.0,1062.5,21.35,4179.1,0,0,95124
1122,0,0,0,0,19,0,No phone service,DSL,0,0,1,1,One year,1,Credit card (automatic),44.85,893.55,1,27,53,0.0,5182,1,San Jose,0,0,Cable,37.294926000000004,-121.89476299999998,0,46.64400000000001,0,0,None,46185,0,0,0,1,19,2,474.0,0.0,0.0,893.55,1,0,95125
1123,1,0,1,1,25,1,0,DSL,1,1,0,0,One year,1,Bank transfer (automatic),61.6,1611,0,46,19,6.45,3807,0,San Jose,1,1,DSL,37.327069,-121.91681899999999,1,61.6,0,5,None,27023,0,0,1,0,25,2,306.0,161.25,44.9,1611.0,0,0,95126
1124,1,0,0,0,12,1,0,DSL,0,1,0,0,Month-to-month,1,Bank transfer (automatic),49.05,593.05,0,58,12,44.78,4244,0,San Jose,0,1,Fiber Optic,37.375156,-121.79586699999999,0,49.05,0,0,None,60620,0,0,0,0,12,3,0.0,537.36,29.32,593.05,0,1,95127
1125,1,1,1,0,39,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.65,4284.8,1,65,29,33.25,4687,1,San Jose,1,1,DSL,37.316146,-121.93628500000001,1,109.876,0,1,None,32804,0,0,1,1,39,4,1243.0,1296.75,0.0,4284.8,0,0,95128
1126,1,0,0,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,74.65,544.55,1,23,78,21.58,3331,1,San Jose,1,1,Cable,37.305622,-122.000887,0,77.63600000000002,0,0,Offer E,37570,0,0,0,1,7,2,425.0,151.06,0.0,544.55,1,0,95129
1127,0,0,1,1,23,1,0,DSL,1,1,0,0,One year,1,Mailed check,66.25,1533.8,0,29,58,11.4,2072,0,San Jose,1,0,DSL,37.277592,-121.98647700000001,1,66.25,0,4,None,13481,1,0,1,0,23,0,890.0,262.2,23.92,1533.8,1,0,95130
1128,1,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.4,529.8,0,26,0,20.66,3792,0,San Jose,0,1,NA,37.387027,-121.897775,0,19.4,0,0,None,26389,0,0,0,0,27,2,0.0,557.82,0.0,529.8,1,0,95131
1129,1,1,0,0,47,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),86.05,3865.6,0,70,20,44.08,5527,0,San Jose,0,1,DSL,37.424655,-121.74841,0,86.05,0,0,None,40568,0,0,0,0,47,1,0.0,2071.76,0.0,3865.6,0,1,95132
1130,1,0,1,1,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.15,515.75,0,45,0,43.84,4347,0,San Jose,0,1,NA,37.371862,-121.860349,1,19.15,2,9,None,26032,0,0,1,0,26,1,0.0,1139.84,0.0,515.75,0,0,95133
1131,0,0,1,0,14,1,1,DSL,1,0,1,0,Month-to-month,1,Bank transfer (automatic),64.7,941,1,51,33,20.4,4049,1,San Jose,0,0,Fiber Optic,37.42765,-121.945416,1,67.28800000000001,0,1,Offer D,9657,0,1,1,0,14,4,0.0,285.6,0.0,941.0,0,1,95134
1132,0,1,1,0,11,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),104.05,1133.65,1,73,30,17.25,4553,1,San Jose,1,0,Cable,37.28682,-121.723877,1,108.212,0,5,None,15798,1,0,1,0,11,1,340.0,189.75,0.0,1133.65,0,0,95135
1133,1,0,0,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.25,48.35,0,58,0,21.18,4725,0,San Jose,0,1,NA,37.270938,-121.851046,0,19.25,1,0,None,36944,0,0,0,0,2,2,0.0,42.36,0.0,48.35,0,0,95136
1134,0,0,1,1,26,1,0,Fiber optic,1,1,0,0,Month-to-month,0,Electronic check,81.95,2070.05,0,23,27,42.95,2817,0,San Jose,0,0,Fiber Optic,37.246064000000004,-121.749494,1,81.95,3,10,None,14792,0,1,1,0,26,1,559.0,1116.7,0.0,2070.05,1,0,95138
1135,0,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.65,8333.95,0,73,27,4.59,5408,0,San Jose,1,0,Fiber Optic,37.218705,-121.762429,1,114.65,0,1,Offer A,7023,1,0,1,0,72,0,2250.0,330.48,0.0,8333.95,0,0,95139
1136,0,0,1,1,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.0,1209.25,0,40,0,46.9,5975,0,Mount Hamilton,0,0,NA,37.382909000000005,-121.634151,1,20.0,2,7,Offer B,38,0,0,1,0,63,1,0.0,2954.7,0.0,1209.25,0,0,95140
1137,1,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.8,1396.25,0,52,0,23.34,5406,0,San Jose,0,1,NA,37.339533,-121.777179,1,19.8,2,9,Offer A,44103,0,0,1,0,71,2,0.0,1657.14,0.0,1396.25,0,0,95148
1138,1,0,1,1,11,1,1,DSL,1,0,1,0,Month-to-month,1,Bank transfer (automatic),65.15,723.35,0,19,59,16.71,5942,0,Stockton,0,1,Fiber Optic,37.959706,-121.287669,1,65.15,2,7,None,7071,0,0,1,0,11,2,42.68,183.81,0.0,723.35,1,1,95202
1139,1,1,1,0,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.65,228.65,0,73,0,45.76,2962,0,Stockton,0,1,NA,37.954089,-121.329761,1,19.65,0,8,None,16357,0,0,1,0,14,0,0.0,640.64,0.0,228.65,0,0,95203
1140,0,0,0,1,13,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),88.95,1161.75,0,30,52,37.03,5407,0,Stockton,1,0,Fiber Optic,37.974498,-121.31956799999999,0,88.95,0,0,None,30476,1,0,0,1,13,2,0.0,481.39,0.0,1161.75,0,1,95204
1141,1,0,0,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.2,98.35,0,38,0,16.91,3478,0,Stockton,0,1,NA,37.965695000000004,-121.260051,0,20.2,2,0,None,34138,0,0,0,0,6,0,0.0,101.46,0.0,98.35,0,0,95205
1142,1,1,1,1,11,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.2,775.3,0,65,22,28.64,5193,0,Stockton,0,1,DSL,37.902421999999994,-121.44002900000001,1,75.2,1,8,None,49657,0,0,1,0,11,0,171.0,315.04,0.0,775.3,0,0,95206
1143,1,0,1,0,18,1,1,DSL,0,1,0,0,Month-to-month,0,Credit card (automatic),56.8,1074.65,0,19,30,1.28,5558,0,Stockton,0,1,Fiber Optic,38.002125,-121.324979,1,56.8,0,5,None,49965,0,0,1,0,18,0,322.0,23.04,0.0,1074.65,1,0,95207
1144,1,0,0,0,1,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,35.55,35.55,1,38,29,0.0,3958,1,Stockton,0,1,Fiber Optic,38.044523,-121.34804799999999,0,36.972,0,0,None,30814,0,1,0,1,1,2,0.0,0.0,0.0,35.55,0,1,95209
1145,0,0,1,0,32,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),75.5,2324.7,0,21,47,19.3,3131,0,Stockton,0,0,DSL,38.033219,-121.29743300000001,1,75.5,0,6,Offer C,40611,0,0,1,0,32,0,0.0,617.6,0.0,2324.7,1,1,95210
1146,1,0,0,0,29,0,No phone service,DSL,1,0,0,0,One year,0,Mailed check,35.6,1072.6,0,46,8,0.0,3898,0,Stockton,0,1,Cable,38.049457000000004,-121.21653,0,35.6,0,0,Offer C,6951,1,0,0,0,29,0,0.0,0.0,0.0,1072.6,0,1,95212
1147,0,0,0,0,3,1,1,DSL,0,0,1,0,Month-to-month,1,Electronic check,60.25,170.5,0,62,29,20.1,4830,0,Stockton,0,0,Fiber Optic,37.946282000000004,-121.139499,0,60.25,0,0,None,23789,0,1,0,0,3,3,0.0,60.3,0.0,170.5,0,1,95215
1148,0,0,0,0,2,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.15,196.9,1,32,28,38.51,2414,1,Stockton,0,0,Fiber Optic,38.029728999999996,-121.387999,0,98.956,0,0,Offer E,19109,0,0,0,1,2,3,55.0,77.02,0.0,196.9,0,0,95219
1149,1,0,1,1,13,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,96.65,1162.85,1,54,12,45.6,5295,1,Acampo,1,1,DSL,38.200231,-121.23503400000001,1,100.516,0,4,Offer D,6317,0,1,1,1,13,1,13.95,592.8000000000002,0.0,1162.85,0,1,95220
1150,0,0,0,0,41,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Electronic check,40.35,1677.85,0,59,21,0.0,2454,0,Angels Camp,0,0,Fiber Optic,38.071327000000004,-120.632221,0,40.35,0,0,Offer B,4264,0,2,0,1,41,1,352.0,0.0,0.0,1677.85,0,0,95222
1151,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,18.85,18.85,0,59,0,7.8,5084,0,Arnold,0,0,NA,38.321529999999996,-120.23635800000001,0,18.85,0,0,None,5159,0,0,0,0,1,0,0.0,7.8,0.0,18.85,0,0,95223
1152,1,0,0,0,7,1,0,DSL,0,0,1,0,Month-to-month,0,Mailed check,54.85,370.4,0,57,24,5.61,3481,0,Avery,0,1,Fiber Optic,38.208335999999996,-120.33993799999999,0,54.85,0,0,None,115,0,0,0,0,7,0,89.0,39.27,0.0,370.4,0,0,95224
1153,0,0,1,0,52,1,0,DSL,1,0,1,0,One year,1,Mailed check,64.3,3410.6,0,36,18,4.22,4405,0,Burson,1,0,Cable,38.183918,-120.898817,1,64.3,0,0,Offer B,27,0,0,0,0,52,3,61.39,219.44,0.0,3410.6,0,1,95225
1154,0,0,1,1,45,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.65,1138.8,0,48,0,20.11,3043,0,Campo Seco,0,0,NA,38.233878999999995,-120.86166599999999,1,24.65,1,7,Offer B,75,0,0,1,0,45,1,0.0,904.95,0.0,1138.8,0,0,95226
1155,1,0,1,0,70,1,1,DSL,0,1,1,0,Two year,0,Credit card (automatic),76.1,5264.25,0,55,9,33.37,5115,0,Clements,1,1,Cable,38.227284999999995,-121.02788999999999,1,76.1,0,4,Offer A,722,1,0,1,0,70,0,474.0,2335.9,0.0,5264.25,0,0,95227
1156,0,0,0,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,18.7,1005.7,0,62,0,10.32,4116,0,Copperopolis,0,0,NA,37.943954,-120.67108,0,18.7,0,0,Offer B,2633,0,0,0,0,53,2,0.0,546.96,0.0,1005.7,0,0,95228
1157,0,1,1,0,62,1,1,Fiber optic,0,1,1,0,One year,1,Credit card (automatic),97.95,5936.55,0,65,25,11.41,5428,0,Farmington,1,0,Fiber Optic,37.956963,-120.863055,1,97.95,0,5,None,596,0,0,1,0,62,0,0.0,707.42,0.0,5936.55,0,1,95230
1158,0,0,1,0,60,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Credit card (automatic),94.1,5475.9,0,44,19,15.54,5267,0,French Camp,0,0,Fiber Optic,37.873283,-121.29203400000002,1,94.1,0,8,Offer B,5094,0,0,1,1,60,1,1040.0,932.4,0.0,5475.9,0,0,95231
1159,0,1,1,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.4,224.05,1,74,10,3.29,3834,1,Glencoe,0,0,Cable,38.358464,-120.57930400000001,1,83.61600000000001,0,1,Offer E,21,0,0,1,0,3,0,0.0,9.87,0.0,224.05,0,1,95232
1160,0,1,1,0,23,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,95.1,2326.05,0,67,12,41.88,4025,0,Hathaway Pines,0,0,Fiber Optic,38.184914,-120.364085,1,95.1,0,1,None,335,0,0,1,1,23,0,279.0,963.24,0.0,2326.05,0,0,95233
1161,1,0,0,1,1,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Mailed check,31.35,31.35,1,41,7,0.0,3605,1,Linden,0,1,DSL,38.047746000000004,-121.030499,0,32.604,0,0,Offer E,3148,0,0,0,0,1,2,0.0,0.0,0.0,31.35,0,0,95236
1162,0,0,0,0,67,1,0,DSL,1,0,0,1,One year,1,Bank transfer (automatic),72.35,4991.5,0,63,9,5.39,4910,0,Lockeford,1,0,DSL,38.166790999999996,-121.14206999999999,0,72.35,0,0,None,3205,1,0,0,1,67,0,0.0,361.13,0.0,4991.5,0,1,95237
1163,0,0,0,0,12,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),89.75,1052.4,1,57,7,14.38,5671,1,Lodi,0,0,Cable,38.123544,-121.15907800000001,0,93.34,0,0,Offer D,45755,0,0,0,0,12,4,74.0,172.56,0.0,1052.4,0,0,95240
1164,0,1,1,0,71,1,1,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),82.7,5831.2,0,72,24,37.53,5089,0,Lodi,1,0,DSL,38.128087,-121.4078,1,82.7,0,1,Offer A,22073,1,0,1,1,71,3,1399.0,2664.63,0.0,5831.2,0,0,95242
1165,1,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.9,510.8,0,41,0,7.17,2130,0,Mokelumne Hill,0,1,NA,38.304194,-120.592431,0,19.9,0,0,Offer C,2718,0,0,0,0,25,2,0.0,179.25,0.0,510.8,0,0,95245
1166,0,0,0,0,5,1,1,DSL,1,0,0,0,Month-to-month,1,Electronic check,53.8,283.95,0,56,22,49.4,2182,0,Mountain Ranch,0,0,Fiber Optic,38.264262,-120.515133,0,53.8,0,0,None,1692,0,0,0,0,5,0,62.0,247.0,0.0,283.95,0,0,95246
1167,1,0,0,0,26,1,1,DSL,0,0,0,0,One year,1,Credit card (automatic),51.55,1295.4,0,29,59,24.67,3130,0,Murphys,0,1,DSL,38.147852,-120.440124,0,51.55,0,0,Offer C,4353,0,0,0,0,26,1,0.0,641.4200000000002,0.0,1295.4,1,1,95247
1168,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.65,19.65,0,21,0,23.41,2539,0,San Andreas,0,1,NA,38.196496999999994,-120.61688999999998,1,19.65,0,1,Offer E,3930,0,1,1,0,1,1,0.0,23.41,0.0,19.65,1,0,95249
1169,1,1,0,0,70,0,No phone service,DSL,0,1,1,0,One year,1,Credit card (automatic),44.05,3011.65,0,68,13,0.0,4022,0,Sheep Ranch,1,1,Fiber Optic,38.244806,-120.417301,0,44.05,0,0,Offer A,88,0,0,0,0,70,2,0.0,0.0,0.0,3011.65,0,1,95250
1170,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,114.0,8093.15,0,60,76,32.47,4558,0,Vallecito,1,1,Fiber Optic,38.055562,-120.456298,1,114.0,3,1,None,460,1,0,1,1,72,0,0.0,2337.84,0.0,8093.15,0,1,95251
1171,1,0,1,0,60,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,94.4,5610.25,1,33,32,47.4,4990,1,Valley Springs,0,1,DSL,38.156971,-120.849231,1,98.17600000000002,0,9,Offer B,11266,0,0,1,1,60,4,0.0,2844.0,0.0,5610.25,0,1,95252
1172,0,1,1,1,32,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.4,3217.65,0,77,19,49.21,4848,0,Wallace,0,0,Fiber Optic,38.192608,-120.957842,1,100.4,2,1,Offer C,304,0,0,1,0,32,1,0.0,1574.72,0.0,3217.65,0,1,95254
1173,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.85,19.85,1,32,0,31.77,3874,1,West Point,0,1,NA,38.41935,-120.469545,0,19.85,0,0,Offer E,2198,0,0,0,0,1,6,0.0,31.77,0.0,19.85,0,0,95255
1174,0,0,0,0,14,1,1,DSL,0,1,0,0,One year,1,Mailed check,54.25,773.2,0,33,7,21.03,4423,0,Wilseyville,0,0,Fiber Optic,38.392686,-120.415951,0,54.25,0,0,Offer D,435,0,0,0,0,14,1,0.0,294.42,0.0,773.2,0,1,95257
1175,0,0,0,0,13,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),80.0,1029.35,0,59,15,33.69,5577,0,Woodbridge,0,0,DSL,38.169605,-121.31096399999998,0,80.0,0,0,Offer D,4176,0,0,0,0,13,2,0.0,437.97,0.0,1029.35,0,1,95258
1176,0,0,0,0,6,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),109.9,669.45,1,55,11,20.36,5750,1,Atwater,1,0,Fiber Optic,37.321233,-120.65635400000001,0,114.296,0,0,Offer E,27808,1,1,0,1,6,3,74.0,122.16,0.0,669.45,0,0,95301
1177,0,0,0,0,46,1,1,DSL,1,0,1,1,Two year,0,Mailed check,79.2,3593.8,0,56,2,46.83,2007,0,Ballico,1,0,Fiber Optic,37.4695,-120.672724,0,79.2,0,0,Offer B,809,0,0,0,1,46,1,7.19,2154.18,0.0,3593.8,0,1,95303
1178,1,0,0,0,15,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.35,1553.95,1,42,13,45.92,3025,1,Big Oak Flat,1,1,Cable,37.818589,-120.25699499999999,0,105.404,0,0,Offer D,167,1,1,0,1,15,2,0.0,688.8000000000002,0.0,1553.95,0,1,95305
1179,1,1,1,0,43,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,94.3,3953.15,0,71,5,4.59,2040,0,Catheys Valley,0,1,Fiber Optic,37.394411,-120.12726200000002,1,94.3,0,1,None,986,1,0,1,0,43,2,198.0,197.37,0.0,3953.15,0,0,95306
1180,1,0,0,0,39,1,0,DSL,0,0,0,0,Two year,1,Bank transfer (automatic),49.8,1971.15,0,59,15,3.93,2202,0,Ceres,0,1,Fiber Optic,37.553469,-120.952825,0,49.8,0,0,Offer C,32881,1,0,0,0,39,0,0.0,153.27,0.0,1971.15,0,1,95307
1181,1,1,0,0,21,1,0,DSL,0,0,1,0,Month-to-month,1,Bank transfer (automatic),60.05,1236.15,1,80,15,34.62,4716,1,Columbia,1,1,Cable,38.085839,-120.37855,0,62.452,0,0,None,2144,0,1,0,0,21,1,185.0,727.02,0.0,1236.15,0,0,95310
1182,1,0,0,0,57,0,No phone service,DSL,1,0,1,1,Month-to-month,1,Electronic check,53.75,3196,0,56,30,0.0,5594,0,Coulterville,1,1,Fiber Optic,37.722127,-120.110174,0,53.75,0,0,Offer B,2271,0,0,0,1,57,0,0.0,0.0,0.0,3196.0,0,1,95311
1183,0,0,1,0,53,1,0,Fiber optic,0,0,1,1,One year,1,Electronic check,93.45,4872.2,0,29,82,38.35,4700,0,Cressey,0,0,Fiber Optic,37.420273,-120.66526999999999,1,93.45,0,1,Offer B,55,1,0,1,1,53,1,3995.0,2032.55,0.0,4872.2,1,0,95312
1184,1,0,1,1,18,1,0,Fiber optic,1,0,1,0,Month-to-month,1,Mailed check,87.9,1500.5,0,32,19,24.16,5192,0,Crows Landing,1,1,DSL,37.435664,-121.04905600000001,1,87.9,1,1,Offer D,1508,0,0,1,0,18,0,0.0,434.88,0.0,1500.5,0,1,95313
1185,0,0,0,0,1,1,1,DSL,0,0,0,1,Month-to-month,1,Electronic check,60.15,60.15,1,19,65,33.48,4611,1,Delhi,0,0,Cable,37.422961,-120.76549299999999,0,62.556000000000004,0,0,Offer E,10159,0,0,0,1,1,5,0.0,33.48,0.0,60.15,1,0,95315
1186,0,0,1,0,58,1,1,DSL,1,0,0,0,One year,1,Bank transfer (automatic),61.05,3478.75,0,59,8,26.36,4411,0,Denair,0,0,Fiber Optic,37.524721,-120.757977,1,61.05,0,1,Offer B,5513,1,0,1,0,58,1,27.83,1528.88,0.0,3478.75,0,1,95316
1187,0,1,0,0,71,1,1,Fiber optic,0,0,1,1,Two year,0,Bank transfer (automatic),104.05,7413.55,0,75,16,47.86,4113,0,El Nido,1,0,Fiber Optic,37.127386,-120.506422,0,104.05,0,0,Offer A,808,0,0,0,0,71,0,1186.0,3398.06,0.0,7413.55,0,0,95317
1188,0,0,0,0,35,1,0,Fiber optic,0,0,1,1,One year,1,Electronic check,99.25,3532,0,38,2,36.42,3244,0,El Portal,1,0,Fiber Optic,37.654551,-119.822984,0,99.25,0,0,Offer C,579,1,0,0,1,35,0,0.0,1274.7,0.0,3532.0,0,1,95318
1189,1,0,0,0,3,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Credit card (automatic),85.7,256.75,0,21,30,29.84,5806,0,Escalon,1,1,Fiber Optic,37.818543,-121.00690700000001,0,85.7,0,0,Offer E,11474,0,0,0,1,3,0,0.0,89.52,0.0,256.75,1,1,95320
1190,1,0,0,0,38,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,104.85,3887.25,0,47,26,4.34,2709,0,Groveland,0,1,Fiber Optic,37.902968,-119.66754399999999,0,104.85,0,0,Offer C,3680,0,0,0,1,38,0,1011.0,164.92,0.0,3887.25,0,0,95321
1191,1,0,1,1,35,1,1,DSL,1,1,0,0,Two year,1,Credit card (automatic),69.15,2490.15,0,60,20,5.06,3945,0,Gustine,1,1,Fiber Optic,37.147197999999996,-121.12016100000001,1,69.15,0,0,Offer C,7872,1,0,0,0,35,0,0.0,177.1,0.0,2490.15,0,1,95322
1192,1,0,0,0,7,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,90.45,593.45,1,31,30,35.91,5356,1,Hickman,1,1,Fiber Optic,37.605926000000004,-120.69955,0,94.068,0,0,Offer E,1055,0,0,0,0,7,4,17.8,251.37,0.0,593.45,0,1,95323
1193,0,0,0,0,47,1,0,DSL,0,0,1,1,Two year,0,Mailed check,74.45,3510.3,0,33,12,3.47,3459,0,Hilmar,1,0,Cable,37.394535999999995,-120.89074699999999,0,74.45,0,0,Offer B,7177,1,1,0,1,47,2,421.0,163.09,0.0,3510.3,0,0,95324
1194,0,0,0,0,14,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,50.45,765.45,0,25,48,39.22,3185,0,Hornitos,0,0,DSL,37.479926,-120.230424,0,50.45,0,0,Offer D,128,0,2,0,0,14,2,0.0,549.0799999999998,0.0,765.45,1,1,95325
1195,0,1,1,0,20,1,0,DSL,0,1,0,1,Month-to-month,1,Electronic check,60.0,1259.35,0,70,16,8.98,2399,0,Hughson,0,0,DSL,37.5923,-120.85328799999999,1,60.0,0,1,None,6822,0,0,1,0,20,0,0.0,179.60000000000005,0.0,1259.35,0,1,95326
1196,1,0,1,0,66,1,1,DSL,1,1,1,1,Two year,0,Electronic check,85.25,5538.35,0,58,21,42.85,5012,0,Jamestown,0,1,DSL,37.84771,-120.486589,1,85.25,0,1,None,9559,1,0,1,1,66,0,0.0,2828.1,0.0,5538.35,0,1,95327
1197,1,0,1,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.45,340.85,0,26,0,39.84,2483,0,Keyes,0,1,NA,37.555631,-120.911653,1,19.45,0,1,Offer D,2130,0,1,1,0,15,2,0.0,597.6,0.0,340.85,1,0,95328
1198,0,0,0,0,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.75,844.45,0,24,0,18.31,2574,0,La Grange,0,0,NA,37.666587,-120.41151699999999,0,20.75,0,0,Offer B,1749,0,0,0,0,42,0,0.0,769.02,0.0,844.45,1,0,95329
1199,0,0,1,0,17,1,1,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,78.9,1348.95,0,53,4,21.15,2362,0,Lathrop,0,0,DSL,37.808209999999995,-121.308401,1,78.9,0,1,Offer D,10834,0,0,1,0,17,0,0.0,359.5499999999999,0.0,1348.95,0,1,95330
1200,1,0,0,0,37,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),104.5,3778,0,26,59,38.72,4812,0,Le Grand,0,1,Cable,37.249377,-120.249581,0,104.5,0,0,Offer C,3256,1,0,0,1,37,0,2229.0,1432.64,0.0,3778.0,1,0,95333
1201,0,0,0,0,12,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,49.4,611.65,0,20,48,17.14,5007,0,Livingston,0,0,Fiber Optic,37.361987,-120.74839399999999,0,49.4,0,0,Offer D,12672,0,0,0,0,12,0,0.0,205.68,0.0,611.65,1,1,95334
1202,1,0,1,0,53,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),94.25,4867.95,1,48,10,15.77,5414,1,Long Barn,0,1,Cable,38.109125,-120.078597,1,98.02,0,1,Offer B,683,0,1,1,1,53,1,487.0,835.81,0.0,4867.95,0,0,95335
1203,0,0,0,0,60,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.0,1505.05,0,63,0,39.41,6355,0,Manteca,0,0,NA,37.830267,-121.20101799999999,0,25.0,0,0,Offer B,36738,0,0,0,0,60,0,0.0,2364.6,0.0,1505.05,0,0,95336
1204,1,0,1,1,18,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),25.55,467.85,0,26,52,0.0,4134,0,Manteca,0,1,Cable,37.750822,-121.238423,1,25.55,2,9,Offer D,19867,0,0,1,0,18,1,243.0,0.0,0.0,467.85,1,0,95337
1205,1,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.9,74.9,1,26,84,1.84,2548,1,Mariposa,0,1,Fiber Optic,37.526790999999996,-119.99436999999999,0,77.89600000000002,0,0,Offer E,10226,0,1,0,1,1,4,0.0,1.84,0.0,74.9,1,0,95338
1206,0,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.15,194.2,0,56,15,5.63,2228,0,Merced,0,0,DSL,37.255637,-120.49353700000002,0,70.15,0,0,None,59289,0,0,0,0,3,1,0.0,16.89,0.0,194.2,0,1,95340
1207,0,0,0,1,9,1,0,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),69.4,571.45,0,23,73,16.77,5108,0,Midpines,0,0,Fiber Optic,37.581496,-119.97276200000002,0,69.4,3,0,Offer E,433,1,0,0,1,9,1,41.72,150.93,0.0,571.45,1,1,95345
1208,0,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.25,80.25,1,34,3,32.92,2502,1,Mi Wuk Village,0,0,Cable,38.121601,-120.13391499999999,0,83.46000000000002,0,0,Offer E,1278,0,0,0,0,1,4,0.0,32.92,0.0,80.25,0,0,95346
1209,1,0,1,0,56,1,1,Fiber optic,1,1,0,0,One year,1,Electronic check,93.15,5253.95,0,45,9,40.33,4778,0,Merced,1,1,Fiber Optic,37.40122,-120.514191,1,93.15,0,1,Offer B,23100,0,0,1,0,56,0,47.29,2258.48,0.0,5253.95,0,1,95348
1210,1,0,1,1,17,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.0,1149.65,1,58,12,44.97,3368,1,Modesto,0,1,Fiber Optic,37.671806,-121.007575,1,71.76,0,1,Offer D,52872,0,0,1,0,17,0,0.0,764.49,0.0,1149.65,0,1,95350
1211,0,0,1,1,11,1,1,DSL,0,0,0,1,Month-to-month,1,Electronic check,66.35,740.8,1,62,13,15.69,2860,1,Modesto,0,0,DSL,37.621458000000004,-121.012295,1,69.00399999999999,0,1,Offer D,47536,1,3,1,1,11,4,96.0,172.59,0.0,740.8,0,0,95351
1212,1,0,0,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.55,521.35,0,25,52,8.95,4704,0,Modesto,0,1,Cable,37.639029,-120.964772,0,69.55,0,0,Offer E,27135,0,1,0,0,7,1,0.0,62.64999999999999,0.0,521.35,1,1,95354
1213,0,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.2,1412.65,0,28,0,42.49,5267,0,Modesto,0,0,NA,37.672906,-120.94659399999999,1,20.2,2,5,None,47613,0,2,1,0,69,1,0.0,2931.81,0.0,1412.65,1,0,95355
1214,1,0,0,0,19,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),86.0,1532.45,1,58,12,20.41,4857,1,Modesto,0,1,Cable,37.716186,-121.02583600000001,0,89.44,0,0,Offer D,26055,0,3,0,1,19,2,184.0,387.79,0.0,1532.45,0,0,95356
1215,0,0,1,1,3,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.3,250.05,1,37,15,48.38,3212,1,Modesto,0,0,Fiber Optic,37.670526,-120.877572,1,83.512,0,1,Offer E,13343,0,0,1,1,3,1,38.0,145.14,0.0,250.05,0,0,95357
1216,1,0,1,1,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.4,1090.6,0,42,0,19.7,6393,0,Modesto,0,1,NA,37.612612,-121.10856799999999,1,20.4,3,3,None,30668,0,0,1,0,54,1,0.0,1063.8,0.0,1090.6,0,0,95358
1217,1,0,1,0,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),23.75,1446.8,0,26,0,32.28,4811,0,Newman,0,1,NA,37.343846,-121.039391,1,23.75,0,6,None,8504,0,0,1,0,62,1,0.0,2001.36,0.0,1446.8,1,0,95360
1218,1,0,0,0,24,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),90.55,2282.55,1,40,6,35.93,5927,1,Oakdale,0,1,Cable,37.785033,-120.776141,0,94.17200000000001,0,0,None,25384,0,0,0,0,24,1,13.7,862.3199999999998,0.0,2282.55,0,1,95361
1219,0,0,1,1,62,1,1,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),70.45,4300.45,0,25,41,36.54,5057,0,Patterson,0,0,DSL,37.410236,-121.32033700000001,1,70.45,3,9,None,15536,0,0,1,1,62,0,1763.0,2265.48,0.0,4300.45,1,0,95363
1220,1,0,0,0,17,1,1,DSL,1,0,0,1,Month-to-month,0,Bank transfer (automatic),65.75,1111.2,0,47,5,47.45,3921,0,Pinecrest,0,1,DSL,38.224869,-119.755729,0,65.75,0,0,Offer D,235,0,0,0,1,17,0,0.0,806.6500000000002,0.0,1111.2,0,1,95364
1221,1,0,0,0,9,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,24.6,190.1,0,24,52,0.0,2323,0,Planada,0,1,Fiber Optic,37.329725,-120.306399,0,24.6,0,0,Offer E,4150,0,0,0,0,9,0,0.0,0.0,0.0,190.1,1,1,95365
1222,1,0,1,1,64,1,0,DSL,1,0,1,0,Two year,0,Mailed check,69.25,4447.75,0,30,51,25.74,4226,0,Ripon,1,1,Fiber Optic,37.750778000000004,-121.13238,1,69.25,0,4,None,12646,1,1,1,0,64,1,0.0,1647.36,0.0,4447.75,0,1,95366
1223,0,0,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.9,143.35,1,30,57,26.87,2101,1,Riverbank,0,0,Cable,37.734971,-120.95427099999999,0,78.936,0,0,None,16525,0,1,0,0,2,1,0.0,53.74,0.0,143.35,0,1,95367
1224,1,0,1,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.85,45.85,1,47,7,14.9,3706,1,Salida,0,1,Fiber Optic,37.713152,-121.08738999999998,1,47.68400000000001,0,1,None,12466,0,0,1,0,1,1,0.0,14.9,0.0,45.85,0,0,95368
1225,0,0,1,0,16,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,49.95,810.2,1,36,32,0.0,4840,1,Snelling,0,0,Fiber Optic,37.521708000000004,-120.42684299999999,1,51.94800000000001,0,1,Offer D,1158,1,0,1,1,16,2,259.0,0.0,0.0,810.2,0,0,95369
1226,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.65,1830.05,0,64,0,24.42,5065,0,Sonora,0,0,NA,37.982715999999996,-120.343732,1,24.65,0,3,None,25340,0,0,1,0,72,0,0.0,1758.2400000000002,0.0,1830.05,0,0,95370
1227,1,0,0,0,30,1,1,Fiber optic,1,1,0,0,One year,0,Bank transfer (automatic),90.4,2820.65,0,62,18,7.19,3171,0,Soulsbyville,1,1,DSL,37.990574,-120.261821,0,90.4,0,0,Offer C,1519,0,0,0,0,30,1,50.77,215.7,0.0,2820.65,0,1,95372
1228,0,0,1,0,49,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Mailed check,100.85,4847.35,0,56,10,44.81,5417,0,Stevinson,0,0,Cable,37.316807,-120.855753,1,100.85,0,3,None,1960,0,0,1,1,49,1,0.0,2195.69,0.0,4847.35,0,1,95374
1229,1,0,1,0,61,1,1,DSL,1,0,0,1,Two year,0,Credit card (automatic),75.35,4729.3,0,21,52,28.8,6466,0,Tracy,1,1,Cable,37.680968,-121.446049,1,75.35,0,10,None,69801,1,0,1,1,61,1,0.0,1756.8,0.0,4729.3,1,1,95376
1230,1,0,1,1,47,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Electronic check,87.2,4017.45,0,54,13,1.09,3760,0,Tuolumne,0,1,Fiber Optic,37.939768,-120.188002,1,87.2,1,7,None,3979,0,0,1,0,47,0,0.0,51.23,0.0,4017.45,0,1,95379
1231,1,0,0,0,20,1,0,DSL,1,0,0,1,Month-to-month,0,Credit card (automatic),64.4,1398.6,0,64,29,12.6,2120,0,Turlock,1,1,DSL,37.474396,-120.87591699999999,0,64.4,0,0,Offer D,40545,0,0,0,1,20,1,0.0,252.0,0.0,1398.6,0,1,95380
1232,1,0,1,1,34,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,78.3,2564.3,1,36,13,13.45,2777,1,Turlock,0,1,Fiber Optic,37.529656,-120.85435700000001,1,81.432,0,1,None,24708,0,0,1,0,34,1,333.0,457.3,0.0,2564.3,0,0,95382
1233,0,0,1,1,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.7,1685.9,0,43,0,30.33,5907,0,Twain Harte,0,0,NA,38.107440999999994,-120.230625,1,24.7,2,8,None,4848,0,0,1,0,70,2,0.0,2123.1,0.0,1685.9,0,0,95383
1234,1,0,0,1,54,1,0,Fiber optic,1,1,1,1,One year,1,Electronic check,105.85,5826.65,0,58,11,20.93,5915,0,Vernalis,0,1,Fiber Optic,37.609095,-121.26338100000001,0,105.85,1,0,None,274,1,0,0,1,54,0,0.0,1130.22,0.0,5826.65,0,1,95385
1235,1,1,1,0,61,1,1,Fiber optic,0,1,1,0,One year,1,Mailed check,98.3,6066.55,0,77,8,2.19,5413,0,Waterford,1,1,Fiber Optic,37.669515999999994,-120.62696399999999,1,98.3,0,2,None,8308,1,0,1,0,61,0,0.0,133.59,0.0,6066.55,0,1,95386
1236,1,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.95,228.4,1,44,25,38.38,4428,1,Escondido,0,1,Cable,33.141265000000004,-116.967221,0,80.028,0,0,None,48690,0,2,0,0,3,2,5.71,115.14,0.0,228.4,0,1,92027
1237,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.45,270.2,0,39,0,22.31,3799,0,Winton,0,1,NA,37.421299,-120.59958700000001,0,19.45,0,0,Offer D,11463,0,0,0,0,13,0,0.0,290.03,0.0,270.2,0,0,95388
1238,0,1,0,0,16,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.15,1529.2,1,76,18,38.75,5913,1,Escondido,0,0,DSL,33.141265000000004,-116.967221,0,99.996,0,0,None,48690,0,0,0,0,16,5,275.0,620.0,0.0,1529.2,0,0,92027
1239,0,0,1,1,3,1,0,DSL,0,1,1,0,Month-to-month,1,Credit card (automatic),58.7,168.6,0,25,51,11.47,3654,0,Santa Rosa,0,0,Fiber Optic,38.460516999999996,-122.79033500000001,1,58.7,2,9,Offer E,36125,0,0,1,0,3,1,0.0,34.410000000000004,0.0,168.6,1,1,95401
1240,1,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.15,536.35,0,43,0,17.64,3848,0,Santa Rosa,0,1,NA,38.488431,-122.752839,0,20.15,0,0,Offer C,40270,0,0,0,0,25,1,0.0,441.0,0.0,536.35,0,0,95403
1241,1,0,0,0,30,1,1,DSL,1,0,0,1,Month-to-month,1,Mailed check,64.5,1888.45,0,58,15,2.64,5039,0,Santa Rosa,0,1,Fiber Optic,38.526941,-122.709096,0,64.5,0,0,None,35057,0,0,0,1,30,0,0.0,79.2,0.0,1888.45,0,1,95404
1242,0,0,1,0,21,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Electronic check,28.5,629.35,0,20,59,0.0,3766,0,Santa Rosa,0,0,DSL,38.439696000000005,-122.66881699999999,1,28.5,0,8,Offer D,22250,0,1,1,0,21,2,37.13,0.0,0.0,629.35,1,1,95405
1243,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.3,45.3,1,49,31,34.37,4568,1,Santa Rosa,0,1,DSL,38.394090999999996,-122.739814,0,47.111999999999995,0,0,None,30876,0,0,0,0,1,7,0.0,34.37,0.0,45.3,0,1,95407
1244,0,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.4,289.3,1,47,0,33.14,5379,1,Santa Rosa,0,0,NA,38.468893,-122.58053899999999,0,19.4,0,0,Offer D,25718,0,0,0,0,15,3,0.0,497.1,0.0,289.3,0,0,95409
1245,1,1,1,0,23,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.45,2117.25,0,76,11,46.82,5272,0,Albion,0,1,Cable,39.225694,-123.717354,1,90.45,0,6,None,1054,0,0,1,0,23,0,0.0,1076.86,0.0,2117.25,0,1,95410
1246,0,0,1,1,45,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,105.15,4730.9,0,63,20,47.48,5915,0,Annapolis,0,0,Cable,38.731055,-123.316553,1,105.15,1,9,None,747,0,1,1,1,45,1,0.0,2136.6,0.0,4730.9,0,1,95412
1247,0,0,1,1,24,1,1,Fiber optic,0,1,0,0,One year,0,Bank transfer (automatic),83.15,2033.05,0,60,53,41.45,2404,0,Boonville,1,0,Fiber Optic,39.025867,-123.38154399999999,1,83.15,3,6,None,1374,0,0,1,0,24,2,0.0,994.8,0.0,2033.05,0,1,95415
1248,0,0,0,0,11,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,90.15,987.95,1,46,3,22.36,5250,1,Branscomb,0,0,Cable,39.710591,-123.682799,0,93.756,0,0,Offer D,176,1,0,0,0,11,0,30.0,245.96,0.0,987.95,0,0,95417
1249,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.05,45.05,1,23,80,48.03,4094,1,Caspar,0,1,Cable,39.361283,-123.784599,0,46.852,0,0,None,333,0,2,0,1,1,2,0.0,48.03,0.0,45.05,1,0,95420
1250,0,0,1,0,56,1,1,Fiber optic,0,0,1,1,Two year,0,Bank transfer (automatic),103.2,5744.35,0,60,13,10.13,4534,0,Cazadero,1,0,DSL,38.578807,-123.19338,1,103.2,0,10,None,1575,1,0,1,1,56,1,74.68,567.2800000000002,0.0,5744.35,0,1,95421
1251,0,0,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,75.8,75.8,1,53,29,14.48,3940,1,Clearlake,0,0,Cable,38.965804,-122.63177900000001,0,78.832,0,0,None,13485,0,3,0,0,1,3,0.0,14.48,0.0,75.8,0,1,95422
1252,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.45,19.45,0,62,0,46.59,5820,0,Clearlake Oaks,0,1,NA,39.07116,-122.598542,0,19.45,0,0,Offer E,3684,0,1,0,0,1,1,0.0,46.59,0.0,19.45,0,0,95423
1253,0,0,0,0,7,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.3,523.15,1,54,18,19.21,3830,1,Cloverdale,0,0,DSL,38.801936,-122.93893500000001,0,82.47200000000001,0,0,None,9210,0,0,0,1,7,0,94.0,134.47,0.0,523.15,0,0,95425
1254,0,1,1,0,55,1,0,Fiber optic,0,0,1,0,Two year,0,Credit card (automatic),88.8,4805.3,0,67,4,33.21,4291,0,Cobb,1,0,Cable,38.838088,-122.73203000000001,1,88.8,0,5,None,1591,1,1,1,0,55,1,192.0,1826.55,0.0,4805.3,0,0,95426
1255,0,0,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,30.9,59.05,1,53,20,0.0,2860,1,Comptche,0,0,Cable,39.239818,-123.565432,0,32.135999999999996,0,0,None,371,1,2,0,0,2,4,12.0,0.0,0.0,59.05,0,0,95427
1256,0,0,1,1,72,1,1,DSL,1,0,1,1,Two year,1,Credit card (automatic),85.9,6110.75,0,39,24,10.87,6361,0,Covelo,1,0,Cable,39.83307,-123.17876499999998,1,85.9,0,9,None,2296,1,0,1,1,72,1,0.0,782.64,0.0,6110.75,0,1,95428
1257,0,1,0,0,45,0,No phone service,DSL,0,0,0,1,One year,0,Electronic check,34.2,1596.6,0,67,4,0.0,5715,0,Dos Rios,0,0,Fiber Optic,39.756049,-123.358701,0,34.2,0,0,Offer B,91,0,1,0,0,45,2,64.0,0.0,0.0,1596.6,0,0,95429
1258,0,0,0,0,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.15,1046.2,0,57,0,3.49,2618,0,Duncans Mills,0,0,NA,38.445603000000006,-123.06375600000001,0,20.15,0,0,None,187,0,0,0,0,47,2,0.0,164.03,0.0,1046.2,0,0,95430
1259,0,1,0,0,46,1,0,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),95.25,4424.2,1,73,33,6.13,3180,1,Lakewood,0,0,Cable,33.840524,-118.148403,0,99.06,0,0,None,30173,0,1,0,0,46,1,1460.0,281.98,0.0,4424.2,0,0,90712
1260,1,0,0,0,2,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,50.3,92.75,0,22,51,18.62,5870,0,Elk,0,1,DSL,39.108252,-123.645121,0,50.3,0,0,Offer E,383,0,0,0,0,2,0,0.0,37.24,0.0,92.75,1,1,95432
1261,0,0,1,0,2,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,80.15,194.55,0,49,23,26.58,5251,0,Forestville,0,0,DSL,38.499302,-122.92443999999999,1,80.15,0,0,Offer E,6216,1,1,0,0,2,1,0.0,53.16,0.0,194.55,0,1,95436
1262,0,0,1,0,12,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,51.25,612.1,0,26,73,46.88,3097,0,Fort Bragg,0,0,Fiber Optic,39.455555,-123.68397900000001,1,51.25,0,1,Offer D,14417,0,1,1,0,12,1,0.0,562.5600000000002,0.0,612.1,1,1,95437
1263,0,1,1,0,68,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),89.6,6127.6,1,70,26,24.13,5651,1,Fulton,0,0,DSL,38.493888,-122.77714099999999,1,93.184,0,1,Offer A,476,0,0,1,0,68,0,0.0,1640.84,0.0,6127.6,0,1,95439
1264,1,0,1,1,69,1,0,Fiber optic,0,0,1,1,Two year,1,Credit card (automatic),95.2,6671.7,0,61,30,12.02,6166,0,Geyserville,0,1,Fiber Optic,38.731771,-123.064272,1,95.2,1,6,None,2349,1,0,1,1,69,0,2002.0,829.38,0.0,6671.7,0,0,95441
1265,1,1,0,1,56,1,0,Fiber optic,1,0,1,1,One year,0,Credit card (automatic),94.8,5264.3,0,71,28,10.57,5693,0,Glen Ellen,0,1,DSL,38.368744,-122.52264199999999,0,94.8,2,0,Offer B,4101,0,0,0,0,56,3,1474.0,591.9200000000002,0.0,5264.3,0,0,95442
1266,0,1,0,0,4,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,80.25,303.7,0,66,4,8.75,3828,0,Glenhaven,0,0,Cable,39.045246,-122.743181,0,80.25,0,0,None,175,0,1,0,0,4,2,12.0,35.0,0.0,303.7,0,0,95443
1267,1,0,1,0,64,1,1,DSL,0,1,1,0,Two year,1,Bank transfer (automatic),76.1,4818.8,0,47,20,6.59,4222,0,Graton,1,1,DSL,38.434362,-122.86891000000001,1,76.1,0,4,None,390,1,0,1,0,64,1,964.0,421.76,0.0,4818.8,0,0,95444
1268,1,0,1,0,59,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,110.15,6448.05,1,43,29,22.71,4601,1,Gualala,1,1,DSL,38.848082,-123.50608000000001,1,114.556,0,1,Offer B,1916,0,3,1,1,59,1,1870.0,1339.89,0.0,6448.05,0,0,95445
1269,1,0,1,1,62,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),115.55,7159.05,0,56,21,40.66,6349,0,Guerneville,1,1,Fiber Optic,38.52576,-123.013347,1,115.55,3,3,None,4913,1,0,1,1,62,0,1503.0,2520.92,0.0,7159.05,0,0,95446
1270,1,0,1,1,63,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.65,1574.5,0,23,0,28.92,4392,0,Healdsburg,0,1,NA,38.618347,-122.908422,1,24.65,2,5,None,17979,0,2,1,0,63,1,0.0,1821.96,0.0,1574.5,1,0,95448
1271,0,0,0,0,53,0,No phone service,DSL,1,1,1,0,One year,1,Electronic check,53.6,2879.2,0,34,25,0.0,5183,0,Hopland,1,0,Fiber Optic,38.937059999999995,-123.11811100000001,0,53.6,0,0,None,1373,1,0,0,0,53,0,720.0,0.0,0.0,2879.2,0,0,95449
1272,1,0,1,1,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.45,86.05,0,20,0,8.04,4573,0,Jenner,0,1,NA,38.505995,-123.18701899999999,1,19.45,1,10,None,438,0,0,1,0,5,0,0.0,40.2,0.0,86.05,1,0,95450
1273,1,1,1,0,49,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,88.2,4159.45,0,75,16,26.0,5987,0,Kelseyville,1,1,DSL,38.93496,-122.792243,1,88.2,0,5,Offer B,9902,0,0,1,0,49,1,0.0,1274.0,0.0,4159.45,0,1,95451
1274,0,0,1,1,62,1,1,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),101.15,6638.35,0,32,52,28.64,5735,0,Kenwood,0,0,Fiber Optic,38.419525,-122.52158500000002,1,101.15,3,4,None,1653,0,0,1,1,62,2,345.19,1775.68,0.0,6638.35,0,1,95452
1275,0,0,1,0,55,1,0,DSL,1,1,0,0,Two year,0,Mailed check,56.8,3112.05,0,28,69,2.36,4702,0,Lakeport,0,0,Fiber Optic,39.080469,-122.955176,1,56.8,0,5,None,11180,1,0,1,0,55,0,2147.0,129.79999999999998,0.0,3112.05,1,0,95453
1276,0,1,1,0,71,1,0,Fiber optic,1,1,1,0,Two year,1,Electronic check,99.4,7168.25,0,78,3,12.26,4964,0,Laytonville,1,0,Cable,39.806141,-123.531098,1,99.4,0,2,Offer A,2706,1,0,1,0,71,0,21.5,870.46,0.0,7168.25,0,1,95454
1277,0,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.1,1326.25,0,25,0,22.05,4603,0,Little River,0,0,NA,39.245911,-123.77214,1,20.1,2,6,None,882,0,0,1,0,72,1,0.0,1587.6,0.0,1326.25,1,0,95456
1278,1,0,1,1,36,0,No phone service,DSL,1,0,1,1,One year,0,Credit card (automatic),60.7,2234.55,0,59,24,0.0,3671,0,Lower Lake,1,1,DSL,38.925545,-122.54908300000001,1,60.7,0,7,None,2644,1,0,1,1,36,1,536.0,0.0,0.0,2234.55,0,0,95457
1279,1,0,1,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.95,495.15,0,47,0,25.08,5682,0,Lucerne,0,1,NA,39.141934,-122.770679,1,20.95,0,3,None,3002,0,1,1,0,25,2,0.0,627.0,0.0,495.15,0,0,95458
1280,0,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.85,8317.95,0,74,25,28.72,4796,0,Manchester,1,0,Cable,38.966713,-123.58641200000001,1,114.85,0,3,Offer A,586,1,0,1,0,72,1,2079.0,2067.84,0.0,8317.95,0,0,95459
1281,0,0,0,0,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.25,679.8,0,44,0,49.85,4904,0,Mendocino,0,0,NA,39.305545,-123.743697,0,19.25,0,0,None,2229,0,0,0,0,36,0,0.0,1794.6,0.0,679.8,0,0,95460
1282,1,0,0,0,1,1,0,DSL,0,0,1,1,Month-to-month,1,Mailed check,62.8,62.8,0,55,29,42.19,2438,0,Middletown,0,1,Fiber Optic,38.787446,-122.58675,0,62.8,0,0,None,7789,0,1,0,1,1,1,0.0,42.19,0.0,62.8,0,0,95461
1283,0,0,1,0,72,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,105.5,7544,0,25,59,21.96,5551,0,Monte Rio,1,0,DSL,38.471049,-123.015549,1,105.5,0,0,None,1537,0,0,0,1,72,1,445.1,1581.12,0.0,7544.0,1,1,95462
1284,1,0,1,1,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.85,1188.25,0,50,0,41.19,6144,0,Navarro,0,1,NA,39.182916,-123.552571,1,19.85,1,2,None,148,0,0,1,0,59,0,0.0,2430.21,0.0,1188.25,0,0,95463
1285,1,1,1,0,7,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.5,676.7,1,75,30,13.63,3077,1,Nice,0,1,Fiber Optic,39.12334,-122.83819799999999,1,93.08,0,1,Offer E,2223,0,2,1,0,7,2,203.0,95.41,0.0,676.7,0,0,95464
1286,0,0,0,0,1,1,0,DSL,0,0,1,1,One year,0,Credit card (automatic),74.1,74.1,0,54,30,36.05,2900,0,Occidental,1,0,Cable,38.415003000000006,-122.998726,0,74.1,0,0,None,1880,1,0,0,1,1,2,0.0,36.05,0.0,74.1,0,0,95465
1287,0,0,1,1,30,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,107.5,3242.5,0,62,18,24.56,3094,0,Philo,1,0,Cable,39.094102,-123.500853,1,107.5,2,9,None,1113,1,0,1,1,30,1,0.0,736.8,0.0,3242.5,0,1,95466
1288,1,0,0,0,64,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.55,1240.15,0,42,0,38.96,6036,0,Point Arena,0,1,NA,38.911299,-123.60958799999999,0,19.55,0,0,None,1352,0,0,0,0,64,1,0.0,2493.44,0.0,1240.15,0,0,95468
1289,1,0,0,0,63,1,1,DSL,1,1,0,0,One year,0,Bank transfer (automatic),68.8,4111.35,0,20,59,38.37,5082,0,Potter Valley,1,1,Cable,39.408634,-123.04551599999999,0,68.8,0,0,None,1884,1,0,0,0,63,0,0.0,2417.31,0.0,4111.35,1,1,95469
1290,1,1,1,0,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),84.45,5899.85,0,75,9,16.72,5856,0,Redwood Valley,1,1,DSL,39.298065,-123.25211000000002,1,84.45,0,3,Offer A,5995,0,0,1,0,72,0,53.1,1203.84,0.0,5899.85,0,1,95470
1291,1,0,1,0,8,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,75.0,632.95,1,20,46,5.34,2587,1,Rio Nido,0,1,Cable,38.522328,-122.97932,1,78.0,0,1,None,298,0,2,1,1,8,1,291.0,42.72,0.0,632.95,1,0,95471
1292,0,0,0,0,62,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),84.5,5193.2,0,60,22,6.05,5466,0,Sebastopol,1,0,Fiber Optic,38.398815,-122.861923,0,84.5,0,0,None,31266,1,0,0,1,62,1,114.25,375.1,0.0,5193.2,0,1,95472
1293,1,0,1,1,67,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),111.2,7530.8,0,19,47,40.96,6060,0,Sonoma,1,1,DSL,38.25485,-122.461799,1,111.2,1,6,None,34314,1,0,1,1,67,2,0.0,2744.32,0.0,7530.8,1,1,95476
1294,1,0,0,0,6,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.75,270.95,1,35,11,41.16,2087,1,Ukiah,0,1,Cable,39.134075,-123.23422,0,46.54,0,0,None,30988,0,2,0,0,6,3,30.0,246.96,0.0,270.95,0,0,95482
1295,0,0,1,1,70,1,1,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),80.6,5460.2,0,37,17,43.81,5880,0,Upper Lake,0,0,DSL,39.220368,-122.907693,1,80.6,0,5,None,2344,1,0,1,1,70,0,0.0,3066.7000000000007,0.0,5460.2,0,1,95485
1296,0,1,0,0,20,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Bank transfer (automatic),80.7,1614.2,0,71,4,21.49,3111,0,Westport,0,0,Fiber Optic,39.724433000000005,-123.767578,0,80.7,0,0,None,309,0,0,0,0,20,2,65.0,429.8,0.0,1614.2,0,0,95488
1297,0,0,0,0,5,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.6,402.5,0,50,25,19.3,3469,0,Willits,0,0,DSL,39.492046,-123.375818,0,75.6,0,0,None,13472,0,0,0,0,5,0,0.0,96.5,0.0,402.5,0,1,95490
1298,0,0,1,1,24,0,No phone service,DSL,1,1,1,1,One year,0,Electronic check,57.6,1367.75,0,42,27,0.0,5623,0,Windsor,1,0,Fiber Optic,38.527297,-122.81004399999999,1,57.6,0,6,None,23701,0,0,1,1,24,2,0.0,0.0,0.0,1367.75,0,1,95492
1299,0,0,1,0,11,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.05,483.7,1,41,33,24.83,3200,1,Witter Springs,0,0,DSL,39.222322999999996,-122.98548799999999,1,45.812,0,1,Offer D,240,0,1,1,0,11,4,160.0,273.13,0.0,483.7,0,0,95493
1300,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),110.6,7962.2,0,55,18,4.32,5444,0,Yorkville,1,1,Fiber Optic,38.888351,-123.23964699999999,1,110.6,0,7,None,335,1,1,1,1,72,1,1433.0,311.04,0.0,7962.2,0,0,95494
1301,0,0,1,1,66,1,0,DSL,1,1,0,0,Two year,1,Credit card (automatic),58.2,3810.8,0,26,59,24.27,5313,0,The Sea Ranch,0,0,DSL,38.696659000000004,-123.43686100000001,1,58.2,0,9,None,752,1,0,1,0,66,1,0.0,1601.82,0.0,3810.8,1,1,95497
1302,0,0,1,1,45,1,0,DSL,1,0,1,1,Two year,1,Mailed check,81.0,3533.6,0,41,29,26.01,2934,0,Eureka,1,0,Fiber Optic,40.796621,-124.15428,1,81.0,0,10,None,23224,1,0,1,1,45,3,1025.0,1170.45,0.0,3533.6,0,0,95501
1303,0,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.7,1396.9,0,47,0,38.39,4131,0,Eureka,0,0,NA,40.737431,-124.108897,1,19.7,3,5,None,23570,0,0,1,0,69,0,0.0,2648.91,0.0,1396.9,0,0,95503
1304,1,1,1,0,15,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),85.6,1345.55,1,74,24,45.25,4981,1,Alderpoint,0,1,DSL,40.166028000000004,-123.584144,1,89.024,0,1,None,261,0,5,1,0,15,3,323.0,678.75,0.0,1345.55,0,0,95511
1305,0,0,0,0,28,1,0,DSL,0,0,1,0,Month-to-month,1,Bank transfer (automatic),59.55,1646.45,0,57,3,38.97,3354,0,Blocksburg,1,0,Fiber Optic,40.309088,-123.668201,0,59.55,0,0,None,199,0,0,0,0,28,1,0.0,1091.16,0.0,1646.45,0,1,95514
1306,0,0,0,0,70,1,1,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),115.55,8127.6,1,30,57,10.21,4838,1,Mckinleyville,1,0,DSL,40.965011,-124.01525500000001,0,120.17200000000001,0,0,Offer A,15921,1,3,0,1,70,2,4633.0,714.7,0.0,8127.6,0,0,95519
1307,0,0,0,0,36,1,0,DSL,1,1,0,1,One year,1,Mailed check,75.55,2680.15,0,48,23,32.0,3235,0,Arcata,1,0,Fiber Optic,40.839958,-124.00375700000001,0,75.55,0,0,None,19596,1,0,0,1,36,1,0.0,1152.0,0.0,2680.15,0,1,95521
1308,1,1,0,0,16,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.6,1281,1,76,24,19.18,2508,1,Bayside,0,1,Cable,40.825486,-124.049485,0,90.064,0,0,None,1689,0,2,0,0,16,2,0.0,306.88,0.0,1281.0,0,1,95524
1309,0,0,0,0,18,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.2,1553.9,1,27,78,24.4,3326,1,Blue Lake,0,0,DSL,40.94338,-123.831799,0,88.60799999999999,0,0,None,1584,0,0,0,1,18,0,0.0,439.2,0.0,1553.9,1,1,95525
1310,0,0,1,0,34,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,97.65,3207.55,1,35,18,43.33,3979,1,Bridgeville,0,0,Cable,40.372532,-123.525626,1,101.556,0,1,None,695,0,0,1,1,34,0,57.74,1473.22,0.0,3207.55,0,1,95526
1311,1,0,1,1,42,0,No phone service,DSL,0,1,0,1,One year,1,Credit card (automatic),45.1,2049.05,0,32,26,0.0,3844,0,Burnt Ranch,1,1,Fiber Optic,40.854512,-123.450097,1,45.1,0,6,None,485,0,0,1,1,42,1,53.28,0.0,0.0,2049.05,0,1,95527
1312,1,0,0,0,48,1,1,DSL,1,0,0,1,One year,1,Bank transfer (automatic),70.95,3629.2,0,50,18,44.76,2667,0,Carlotta,0,1,Fiber Optic,40.497283,-123.93037,0,70.95,0,0,Offer B,1072,1,0,0,1,48,3,0.0,2148.48,0.0,3629.2,0,1,95528
1313,1,0,1,0,47,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,109.55,5124.55,1,54,22,7.62,5863,1,Fallbrook,1,1,DSL,33.362575,-117.299644,1,113.932,0,1,Offer B,42239,1,0,1,1,47,2,1127.0,358.14,0.0,5124.55,0,0,92028
1314,0,0,1,1,39,1,1,Fiber optic,0,1,0,0,One year,1,Electronic check,89.55,3474.45,1,50,33,35.32,3849,1,Ferndale,1,0,Cable,40.4785,-124.301372,1,93.132,0,1,None,2965,1,0,1,0,39,5,1147.0,1377.48,0.0,3474.45,0,0,95536
1315,0,0,1,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.9,202.3,0,32,0,2.52,5359,0,Fields Landing,0,0,NA,40.726949,-124.217378,1,20.9,1,3,Offer D,228,0,0,1,0,11,0,0.0,27.72,0.0,202.3,0,0,95537
1316,1,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.95,147.5,0,47,0,13.86,3331,0,Fortuna,0,1,NA,40.584990999999995,-124.121504,0,19.95,0,0,None,12241,0,0,0,0,7,1,0.0,97.02,0.0,147.5,0,0,95540
1317,0,0,0,0,3,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,24.6,86.35,0,27,0,26.33,5756,0,Garberville,0,0,NA,40.057784000000005,-123.679461,0,24.6,0,0,None,2423,0,0,0,0,3,0,0.0,78.99,0.0,86.35,1,0,95542
1318,1,0,0,0,8,1,0,DSL,1,0,0,1,Month-to-month,1,Electronic check,66.7,579,0,47,27,41.13,4490,0,Gasquet,1,1,Fiber Optic,41.867908,-123.79414399999999,0,66.7,0,0,None,532,0,0,0,1,8,0,0.0,329.04,0.0,579.0,0,1,95543
1319,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.45,19.45,1,42,0,48.96,5687,1,Honeydew,0,1,NA,40.342928,-124.06332900000001,0,19.45,0,0,Offer E,82,0,0,0,0,1,2,0.0,48.96,0.0,19.45,0,0,95545
1320,1,0,1,1,32,1,0,Fiber optic,1,1,0,1,One year,0,Mailed check,94.8,3131.55,0,42,76,43.37,5288,0,Hoopa,1,1,DSL,41.163637,-123.70484099999999,1,94.8,3,1,None,3041,0,0,1,1,32,0,238.0,1387.84,0.0,3131.55,0,1,95546
1321,1,0,1,1,60,1,0,DSL,1,1,0,0,One year,1,Bank transfer (automatic),65.85,3928.3,0,35,30,43.57,4053,0,Hydesville,1,1,Fiber Optic,40.557314,-124.08166200000001,1,65.85,0,4,Offer B,1201,1,0,1,0,60,2,1178.0,2614.2,0.0,3928.3,0,0,95547
1322,0,0,1,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.95,187.75,0,21,0,49.6,3831,0,Klamath,0,0,NA,41.572813000000004,-124.03501100000001,1,19.95,0,9,Offer D,1215,0,0,1,0,10,1,0.0,496.0,0.0,187.75,1,0,95548
1323,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.65,1710.15,0,33,0,43.37,4015,0,Kneeland,0,0,NA,40.664483000000004,-123.865325,1,24.65,0,5,None,264,0,0,1,0,71,1,0.0,3079.27,0.0,1710.15,0,0,95549
1324,0,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,76.35,1,34,0,12.43,4133,1,Korbel,0,0,NA,40.7666,-123.80458,1,20.35,0,0,Offer E,155,0,2,0,0,4,3,0.0,49.72,0.0,76.35,0,0,95550
1325,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.25,69.25,1,75,20,29.68,4371,1,Loleta,0,0,Cable,40.665952000000004,-124.240051,0,72.02,0,0,Offer E,1447,0,1,0,0,1,3,0.0,29.68,0.0,69.25,0,0,95551
1326,0,0,1,1,43,0,No phone service,DSL,1,1,1,0,One year,1,Bank transfer (automatic),51.25,2151.6,0,61,6,0.0,5656,0,Mad River,0,0,DSL,40.390301,-123.412327,1,51.25,0,2,Offer B,265,1,0,1,0,43,1,0.0,0.0,0.0,2151.6,0,1,95552
1327,1,0,1,0,59,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),99.5,5961.1,1,33,6,10.76,6098,1,Miranda,1,1,Cable,40.210895,-123.86,1,103.48,0,1,Offer B,867,0,1,1,1,59,3,358.0,634.84,0.0,5961.1,0,0,95553
1328,0,0,1,0,23,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,54.25,1221.55,0,47,4,38.93,5140,0,Myers Flat,1,0,DSL,40.267158,-123.80591299999999,1,54.25,0,6,Offer D,644,1,0,1,0,23,3,0.0,895.39,0.0,1221.55,0,1,95554
1329,0,0,1,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.4,1496.45,0,28,0,12.87,5398,0,Orick,0,0,NA,41.336354,-124.044354,1,19.4,0,8,None,494,0,0,1,0,72,0,0.0,926.64,0.0,1496.45,1,0,95555
1330,1,0,1,0,22,1,0,DSL,1,0,0,0,One year,1,Credit card (automatic),56.25,1292.2,0,56,7,7.68,3733,0,Orleans,0,1,DSL,41.269521000000005,-123.546958,1,56.25,0,8,Offer D,574,1,0,1,0,22,0,9.05,168.95999999999995,0.0,1292.2,0,1,95556
1331,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,25.15,25.15,0,19,52,0.0,3513,0,Petrolia,0,0,Fiber Optic,40.274302,-124.210902,0,25.15,0,0,None,300,0,0,0,0,1,2,0.0,0.0,0.0,25.15,1,0,95558
1332,1,0,0,0,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),23.95,1713.1,0,57,0,22.24,6059,0,Phillipsville,0,1,NA,40.184094,-123.74548700000001,0,23.95,0,0,None,163,0,0,0,0,69,1,0.0,1534.56,0.0,1713.1,0,0,95559
1333,1,0,0,0,50,0,No phone service,DSL,1,0,0,0,One year,1,Mailed check,35.4,1748.9,0,45,7,0.0,5052,0,Redway,0,1,Fiber Optic,40.142256,-123.85292700000001,0,35.4,0,0,Offer B,1851,1,0,0,0,50,1,0.0,0.0,0.0,1748.9,0,1,95560
1334,0,1,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,25.2,25.2,1,74,6,0.0,5688,1,Rio Dell,0,0,DSL,40.485849,-124.163234,0,26.208000000000002,0,0,None,3284,0,1,0,0,1,2,0.0,0.0,0.0,25.2,0,0,95562
1335,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.0,96.45,1,44,3,17.25,5704,1,Salyer,0,1,Fiber Optic,40.89866,-123.539754,0,46.8,0,0,None,660,0,4,0,0,2,1,3.0,34.5,0.0,96.45,0,0,95563
1336,0,0,1,0,15,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),75.35,1114.55,0,22,71,30.09,4891,0,Samoa,0,0,DSL,40.809636,-124.189977,1,75.35,0,6,None,395,0,0,1,0,15,0,0.0,451.35,0.0,1114.55,1,1,95564
1337,1,0,0,0,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.4,609.1,0,56,0,25.58,5363,0,Scotia,0,1,NA,40.440636,-124.098739,0,20.4,0,0,None,1125,0,0,0,0,31,0,0.0,792.9799999999998,0.0,609.1,0,0,95565
1338,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.15,20.15,1,35,0,40.51,4103,1,Smith River,0,1,NA,41.950683000000005,-124.097094,0,20.15,0,0,Offer E,2020,0,0,0,0,1,2,0.0,40.51,0.0,20.15,0,0,95567
1339,1,0,1,0,66,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),105.0,7133.25,1,28,56,7.28,5723,1,Somes Bar,1,1,Cable,41.444606,-123.47189499999999,1,109.2,0,0,Offer A,202,0,2,0,1,66,3,0.0,480.48,0.0,7133.25,1,1,95568
1340,0,0,1,1,0,0,No phone service,DSL,1,1,1,0,Two year,0,Credit card (automatic),56.05, ,0,64,8,0.0,4740,0,Redcrest,1,0,DSL,40.363446,-123.83504099999999,1,56.05,0,2,None,400,1,0,1,0,10,0,0.0,0.0,0.0,560.5,0,1,95569
1341,1,0,0,1,3,1,0,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),54.7,169.45,1,58,19,2.88,3335,1,Trinidad,0,1,Fiber Optic,41.162295,-124.027381,0,56.88800000000001,0,0,Offer E,2369,0,4,0,0,3,4,3.22,8.64,0.0,169.45,0,1,95570
1342,0,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.0,141.6,0,55,0,23.46,3087,0,Weott,0,0,NA,40.310119,-123.909449,0,20.0,0,0,None,270,0,0,0,0,8,2,0.0,187.68,0.0,141.6,0,0,95571
1343,1,0,1,1,64,1,0,DSL,1,0,1,1,One year,1,Credit card (automatic),73.05,4688.65,0,20,71,26.64,4515,0,Willow Creek,1,1,Fiber Optic,40.949011999999996,-123.655847,1,73.05,0,5,Offer B,1666,0,0,1,1,64,0,0.0,1704.96,0.0,4688.65,1,1,95573
1344,0,0,1,0,28,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.5,563.05,0,27,0,42.33,5145,0,Leggett,0,0,NA,39.873371,-123.741474,1,20.5,0,3,None,321,0,0,1,0,28,1,0.0,1185.24,0.0,563.05,1,0,95585
1345,0,0,1,0,57,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),100.75,5985,0,39,11,3.72,6354,0,Piercy,1,0,Fiber Optic,39.955587,-123.681175,1,100.75,0,5,Offer B,200,0,0,1,1,57,0,65.84,212.04,0.0,5985.0,0,1,95587
1346,0,0,1,1,14,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,87.25,1258.6,1,49,21,29.18,4786,1,Fallbrook,1,0,Fiber Optic,33.362575,-117.299644,1,90.74,0,1,None,42239,0,0,1,1,14,2,264.0,408.52,0.0,1258.6,0,0,92028
1347,1,0,0,0,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.95,373.5,0,58,0,19.1,2831,0,Zenia,0,1,NA,40.170357,-123.417298,0,19.95,0,0,None,259,0,0,0,0,19,0,0.0,362.9,0.0,373.5,0,0,95595
1348,1,0,1,0,10,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.95,857.2,1,38,4,11.3,5640,1,Amador City,0,1,DSL,38.431407,-120.8421,1,83.14800000000002,0,1,None,222,0,1,1,0,10,6,34.0,113.0,0.0,857.2,0,0,95601
1349,0,0,1,0,51,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,49.65,2553.35,0,21,42,0.0,5528,0,Auburn,0,0,Fiber Optic,38.99003,-121.11440800000001,1,49.65,0,0,Offer B,18197,0,0,0,1,51,0,0.0,0.0,0.0,2553.35,1,1,95602
1350,0,0,1,0,67,1,1,DSL,1,1,0,0,Two year,0,Mailed check,65.65,4322.85,0,51,22,22.83,5441,0,Auburn,1,0,DSL,38.912881,-121.08276599999999,1,65.65,0,5,None,24944,0,0,1,0,67,0,0.0,1529.61,0.0,4322.85,0,1,95603
1351,1,0,1,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.45,250.8,0,43,0,16.67,2606,0,West Sacramento,0,1,NA,38.592745,-121.54003600000001,1,20.45,2,3,None,12756,0,0,1,0,11,0,0.0,183.37,0.0,250.8,0,0,95605
1352,1,0,1,1,72,0,No phone service,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),60.95,4549.05,0,38,15,0.0,4147,0,Brooks,1,1,Cable,38.809804,-122.24138300000001,1,60.95,0,8,None,382,1,0,1,1,72,0,682.0,0.0,0.0,4549.05,0,0,95606
1353,1,0,1,1,66,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,20.35,1359.5,0,59,0,45.03,4845,0,Capay,0,1,NA,38.681651,-122.130569,1,20.35,0,9,Offer A,262,0,0,1,0,66,0,0.0,2971.98,0.0,1359.5,0,0,95607
1354,0,0,0,0,18,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,88.35,1639.3,1,47,25,12.67,5727,1,Carmichael,0,0,Cable,38.626128,-121.328011,0,91.884,0,0,None,58830,1,2,0,0,18,3,410.0,228.06,0.0,1639.3,0,0,95608
1355,0,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.5,178.85,0,43,0,46.94,4283,0,Citrus Heights,0,0,NA,38.69508,-121.271616,0,19.5,0,0,None,43718,0,0,0,0,9,1,0.0,422.46,0.0,178.85,0,0,95610
1356,0,0,0,0,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.2,633.85,0,59,28,9.27,5841,0,Clarksburg,0,0,DSL,38.384648,-121.578701,0,75.2,0,0,None,1417,0,0,0,0,9,0,0.0,83.42999999999998,0.0,633.85,0,1,95612
1357,1,0,1,0,48,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),111.45,5315.1,0,28,59,22.36,2319,0,Cool,1,1,Fiber Optic,38.880621999999995,-120.97386499999999,1,111.45,0,9,Offer B,3674,0,0,1,1,48,2,0.0,1073.28,0.0,5315.1,1,1,95614
1358,1,0,0,0,10,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.15,735.5,0,23,85,4.29,3963,0,Courtland,0,1,Fiber Optic,38.311609000000004,-121.554034,0,70.15,0,0,None,699,0,0,0,0,10,1,625.0,42.9,0.0,735.5,1,0,95615
1359,0,0,0,0,9,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.75,889.9,1,34,29,10.07,2893,1,Davis,0,0,Cable,38.508734999999994,-121.67881299999999,0,98.54,0,0,Offer E,67411,0,0,0,1,9,1,0.0,90.63,0.0,889.9,0,1,95616
1360,0,1,0,0,13,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.05,1290,1,73,26,19.03,2230,1,Davis,0,0,DSL,38.544002,-121.68555900000001,0,98.852,0,0,None,648,0,0,0,1,13,3,335.0,247.39,0.0,1290.0,0,0,95618
1361,1,0,0,0,4,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,78.45,330.05,1,28,64,42.06,5048,1,Diamond Springs,0,1,Cable,38.683605,-120.811852,0,81.58800000000002,0,0,Offer E,4426,0,0,0,1,4,1,211.0,168.24,0.0,330.05,1,0,95619
1362,1,0,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.2,237.95,1,43,16,13.02,5094,1,Dixon,0,1,Fiber Optic,38.392821000000005,-121.799917,0,73.00800000000002,0,0,None,18529,0,1,0,0,4,3,38.0,52.08,0.0,237.95,0,0,95620
1363,0,0,1,0,72,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),92.0,6474.4,0,47,16,43.29,6434,0,Citrus Heights,1,0,Fiber Optic,38.69549,-121.307864,1,92.0,0,8,Offer A,41636,1,0,1,1,72,1,0.0,3116.88,0.0,6474.4,0,1,95621
1364,0,0,1,1,51,1,0,DSL,1,1,1,1,Two year,0,Credit card (automatic),85.5,4421.95,0,63,13,33.93,6261,0,El Dorado,1,0,Fiber Optic,38.63153,-120.84260900000001,1,85.5,0,10,Offer B,4097,1,0,1,1,51,1,575.0,1730.43,0.0,4421.95,0,0,95623
1365,1,0,1,0,59,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Bank transfer (automatic),41.05,2452.7,1,23,76,0.0,4324,1,Elk Grove,0,1,Fiber Optic,38.434138,-121.30587,1,42.692,0,1,Offer B,38534,0,0,1,1,59,3,1864.0,0.0,0.0,2452.7,1,0,95624
1366,1,0,1,0,10,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.6,813.85,1,63,32,30.1,5146,1,Elmira,0,1,Fiber Optic,38.349195,-121.902943,1,89.024,0,1,None,171,0,1,1,0,10,6,26.04,301.0,0.0,813.85,0,1,95625
1367,1,1,1,0,61,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,82.15,4904.85,0,66,2,26.55,4250,0,Elverta,0,1,Fiber Optic,38.734997,-121.463719,1,82.15,0,4,Offer B,6197,0,0,1,0,61,0,9.81,1619.55,0.0,4904.85,0,1,95626
1368,1,0,0,0,54,1,0,Fiber optic,1,0,0,0,One year,0,Electronic check,84.4,4484.05,0,41,18,30.66,4154,0,Esparto,1,1,DSL,38.834469,-122.12719299999999,0,84.4,0,0,Offer B,2756,1,0,0,0,54,2,80.71,1655.64,0.0,4484.05,0,1,95627
1369,0,0,0,0,33,1,1,DSL,1,1,0,0,Month-to-month,1,Mailed check,60.9,2033.85,0,38,24,15.69,3009,0,Fair Oaks,0,0,DSL,38.652065,-121.25441000000001,0,60.9,0,0,None,40750,0,0,0,0,33,1,0.0,517.77,0.0,2033.85,0,1,95628
1370,0,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.25,538.2,0,62,0,35.77,5250,0,Fiddletown,0,0,NA,38.513484000000005,-120.704613,0,20.25,0,0,None,850,0,0,0,0,27,2,0.0,965.79,0.0,538.2,0,0,95629
1371,0,1,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.2,79.2,1,69,26,20.06,4363,1,Folsom,0,0,DSL,38.672638,-121.147403,0,82.36800000000002,0,0,None,51855,0,0,0,0,1,2,0.0,20.06,0.0,79.2,0,0,95630
1372,1,0,0,0,23,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Mailed check,95.3,2192.9,0,53,23,48.21,5029,0,Foresthill,0,1,DSL,39.031876000000004,-120.81114099999999,0,95.3,0,0,None,5714,0,0,0,1,23,2,0.0,1108.83,0.0,2192.9,0,1,95631
1373,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,19.85,0,63,0,29.1,4840,0,Galt,0,1,NA,38.274451,-121.259201,0,19.85,2,0,None,24194,0,2,0,0,1,1,0.0,29.1,0.0,19.85,0,0,95632
1374,1,0,1,1,45,1,0,DSL,1,1,1,1,Two year,1,Mailed check,84.35,3858.05,0,63,3,30.8,3403,0,Garden Valley,1,1,DSL,38.852544,-120.83766899999999,1,84.35,0,3,Offer B,2536,1,0,1,1,45,0,0.0,1386.0,0.0,3858.05,0,1,95633
1375,0,0,1,1,39,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.85,854.8,0,35,0,32.57,3032,0,Georgetown,0,0,NA,38.9386,-120.78551399999999,1,19.85,1,3,None,2723,0,0,1,0,39,0,0.0,1270.23,0.0,854.8,0,0,95634
1376,1,0,0,0,5,1,0,DSL,0,0,1,1,One year,1,Mailed check,70.0,347.4,1,39,24,45.25,2673,1,Greenwood,1,1,DSL,38.921333000000004,-120.897718,0,72.8,0,0,None,1140,0,0,0,1,5,0,83.0,226.25,0.0,347.4,0,0,95635
1377,1,0,1,1,72,1,1,DSL,1,1,1,0,Two year,0,Bank transfer (automatic),82.3,5815.15,0,40,15,48.44,4162,0,Grizzly Flats,1,1,Fiber Optic,38.636102,-120.522149,1,82.3,0,10,Offer A,659,1,2,1,0,72,2,872.0,3487.68,0.0,5815.15,0,0,95636
1378,0,0,1,1,58,1,1,DSL,0,1,1,0,Month-to-month,1,Bank transfer (automatic),66.8,3970.4,0,44,19,44.1,6433,0,Guinda,0,0,DSL,38.830739,-122.196202,1,66.8,1,2,Offer B,228,0,0,1,0,58,0,0.0,2557.8,0.0,3970.4,0,1,95637
1379,0,0,0,0,70,0,No phone service,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),44.6,3058.15,0,62,11,0.0,4442,0,Herald,1,0,Cable,38.313447,-121.12388600000001,0,44.6,0,0,Offer A,1745,1,0,0,0,70,1,0.0,0.0,0.0,3058.15,0,1,95638
1380,1,0,1,1,61,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),98.45,6145.2,0,41,21,41.57,4000,0,Hood,0,1,Fiber Optic,38.375325,-121.507935,1,98.45,1,4,Offer B,213,1,0,1,1,61,0,0.0,2535.77,0.0,6145.2,0,1,95639
1381,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.7,129.2,0,37,14,2.72,2388,0,Ione,0,1,DSL,38.33788,-120.954202,0,70.7,0,0,Offer E,9752,0,0,0,0,2,1,0.0,5.44,0.0,129.2,0,1,95640
1382,0,0,1,1,46,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,24.95,1165.9,0,39,0,4.6,3979,0,Isleton,0,0,NA,38.154823,-121.601358,1,24.95,0,0,Offer B,2010,0,0,0,0,46,0,0.0,211.6,0.0,1165.9,0,0,95641
1383,0,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),49.95,49.95,1,51,4,43.49,2041,1,Jackson,0,0,Fiber Optic,38.336216,-120.76901000000001,0,51.94800000000001,0,0,None,6202,0,0,0,0,1,0,0.0,43.49,0.0,49.95,0,0,95642
1384,0,0,1,0,22,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.25,1554,1,19,57,32.11,2159,1,Knights Landing,0,0,Cable,38.875508,-121.76586599999999,1,72.02,0,1,None,1793,0,0,1,0,22,0,886.0,706.42,0.0,1554.0,1,0,95645
1385,0,0,0,0,48,1,0,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),102.5,4904.25,0,43,21,19.04,3262,0,Kirkwood,1,0,Cable,38.631489,-120.01516699999999,0,102.5,0,0,Offer B,129,1,0,0,1,48,1,0.0,913.92,0.0,4904.25,0,1,95646
1386,1,0,0,0,64,1,1,DSL,0,1,1,1,Two year,0,Credit card (automatic),86.55,5632.55,0,35,7,14.39,4934,0,Lincoln,1,1,Fiber Optic,38.922812,-121.312005,0,86.55,0,0,Offer B,15286,1,0,0,1,64,3,394.0,920.96,0.0,5632.55,0,0,95648
1387,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.3,1643.25,0,53,0,20.42,5160,0,Loomis,0,1,NA,38.809175,-121.171375,1,24.3,3,3,Offer A,11191,0,1,1,0,72,2,0.0,1470.2400000000002,0.0,1643.25,0,0,95650
1388,0,0,1,1,12,1,0,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),58.35,740.55,0,51,52,7.97,5068,0,Lotus,1,0,Cable,38.815515000000005,-120.916997,1,58.35,3,2,None,485,0,0,1,0,12,1,0.0,95.64,0.0,740.55,0,1,95651
1389,0,1,1,0,34,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,94.25,3217.55,1,75,4,2.88,3369,1,Madison,1,0,Fiber Optic,38.674276,-121.96186599999999,1,98.02,0,1,None,844,0,2,1,0,34,2,0.0,97.92,0.0,3217.55,0,1,95653
1390,0,0,1,1,72,1,0,DSL,1,1,0,1,Two year,0,Credit card (automatic),68.75,4888.2,0,29,59,12.32,4505,0,Mather,1,0,Cable,38.549822,-121.266725,1,68.75,0,6,Offer A,929,0,0,1,1,72,0,2884.0,887.04,0.0,4888.2,1,0,95655
1391,1,0,1,0,29,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,85.8,2440.25,0,62,16,39.5,2568,0,Newcastle,1,1,Fiber Optic,38.883224,-121.15918,1,85.8,0,4,None,6096,0,0,1,0,29,2,390.0,1145.5,0.0,2440.25,0,0,95658
1392,1,0,1,1,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.1,620.55,0,21,0,49.37,3636,0,Nicolaus,0,1,NA,38.788897999999996,-121.608624,1,20.1,0,3,None,751,0,0,1,0,33,0,0.0,1629.2099999999996,0.0,620.55,1,0,95659
1393,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,20.35,0,47,0,44.09,5774,0,North Highlands,0,0,NA,38.671295,-121.388251,0,20.35,0,0,None,32202,0,0,0,0,1,0,0.0,44.09,0.0,20.35,0,0,95660
1394,0,0,1,1,62,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,110.8,6840.95,0,42,57,13.25,4306,0,Roseville,1,0,DSL,38.736684999999994,-121.25198400000001,1,110.8,3,5,Offer B,25173,1,0,1,1,62,1,3899.0,821.5,0.0,6840.95,0,0,95661
1395,1,0,1,0,41,1,1,DSL,0,0,1,1,One year,1,Electronic check,73.0,3001.2,1,34,32,15.91,2041,1,Orangevale,1,1,Cable,38.689174,-121.21843500000001,1,75.92,0,1,None,32040,0,0,1,1,41,4,0.0,652.3100000000002,0.0,3001.2,0,1,95662
1396,0,0,0,0,64,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),100.05,6254.2,1,39,20,28.13,5452,1,Penryn,1,0,Fiber Optic,38.859093,-121.182872,0,104.052,0,0,None,2048,0,3,0,1,64,7,1251.0,1800.32,0.0,6254.2,0,0,95663
1397,0,0,0,0,4,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),82.85,319.6,0,24,73,19.84,3154,0,Pilot Hill,1,0,Fiber Optic,38.803731,-121.04379899999999,0,82.85,0,0,Offer E,1173,0,0,0,1,4,0,0.0,79.36,0.0,319.6,1,1,95664
1398,0,0,0,0,24,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,84.35,1938.05,0,44,3,25.81,2198,0,Pine Grove,0,0,Cable,38.400264,-120.641274,0,84.35,0,0,None,4354,1,0,0,0,24,0,58.0,619.4399999999998,0.0,1938.05,0,0,95665
1399,0,0,1,1,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.55,294.5,0,56,0,19.03,5620,0,Pioneer,0,0,NA,38.546999,-120.27111399999998,1,19.55,0,9,None,5501,0,0,1,0,14,0,0.0,266.42,0.0,294.5,0,0,95666
1400,1,0,0,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,58.3,0,38,0,5.15,4430,0,Placerville,0,1,NA,38.733714,-120.79521299999999,0,19.95,3,0,Offer E,34146,0,0,0,0,3,0,0.0,15.45,0.0,58.3,0,0,95667
1401,0,1,0,0,4,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),99.8,442.85,1,65,11,12.68,2268,1,Pleasant Grove,1,0,Cable,38.833554,-121.498102,0,103.792,0,0,None,901,0,1,0,1,4,4,49.0,50.72,0.0,442.85,0,0,95668
1402,0,0,0,1,18,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,35.0,553,1,27,94,0.0,2649,1,Plymouth,0,0,Cable,38.489273,-120.89161399999999,0,36.4,0,0,None,2220,0,0,0,1,18,2,520.0,0.0,0.0,553.0,1,0,95669
1403,1,0,0,0,8,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,66.25,546.45,0,40,24,25.72,3026,0,Rancho Cordova,0,1,Fiber Optic,38.602723,-121.279913,0,66.25,0,0,Offer E,49729,0,0,0,1,8,2,131.0,205.76,0.0,546.45,0,0,95670
1404,0,0,0,0,35,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),23.3,797.1,0,38,0,6.52,2416,0,Rescue,0,0,NA,38.724321999999994,-120.99123700000001,0,23.3,0,0,None,3815,0,0,0,0,35,1,0.0,228.2,0.0,797.1,0,0,95672
1405,0,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,76.0,76,1,20,57,35.01,2567,1,Rio Linda,0,0,Cable,38.688764,-121.457596,0,79.04,0,0,None,14010,0,1,0,0,1,3,0.0,35.01,0.0,76.0,1,1,95673
1406,1,0,0,1,66,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.3,1673.8,0,64,0,23.81,6019,0,Rio Oso,0,1,NA,38.954144,-121.48253600000001,0,25.3,3,0,Offer A,947,0,2,0,0,66,1,0.0,1571.4599999999996,0.0,1673.8,0,0,95674
1407,1,0,0,1,8,0,No phone service,DSL,1,0,0,1,Two year,1,Mailed check,44.55,343.45,0,46,4,0.0,5489,0,River Pines,0,1,Fiber Optic,38.545775,-120.743325,0,44.55,0,0,None,364,1,0,0,1,8,1,0.0,0.0,0.0,343.45,0,1,95675
1408,0,0,1,0,71,1,1,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),104.1,7412.25,0,19,82,4.39,4695,0,Rocklin,1,0,Fiber Optic,38.7904,-121.23697299999999,1,104.1,0,8,Offer A,21510,0,0,1,1,71,0,6078.0,311.69,0.0,7412.25,1,0,95677
1409,0,0,1,1,43,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),92.55,4039,0,59,53,27.49,3853,0,Roseville,1,0,DSL,38.759751,-121.288545,1,92.55,3,3,Offer B,30614,0,0,1,1,43,0,0.0,1182.07,0.0,4039.0,0,1,95678
1410,0,1,0,0,2,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.85,170.85,1,77,20,19.27,4193,1,Sheridan,0,0,DSL,38.984756,-121.345074,0,97.604,0,0,None,1219,0,0,0,0,2,4,3.42,38.54,0.0,170.85,0,1,95681
1411,1,1,0,0,29,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),101.45,2948.6,0,79,21,6.59,5285,0,Shingle Springs,1,1,Fiber Optic,38.598936,-120.96309199999999,0,101.45,0,0,Offer C,24738,0,0,0,0,29,0,0.0,191.11,0.0,2948.6,0,1,95682
1412,0,0,1,0,15,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.3,1308.4,1,36,31,28.3,4003,1,Sloughhouse,1,0,DSL,38.470423,-121.114897,1,87.67200000000001,0,1,None,4731,0,0,1,0,15,0,0.0,424.5,0.0,1308.4,0,1,95683
1413,1,0,1,1,65,1,1,Fiber optic,1,1,0,0,Two year,0,Credit card (automatic),94.55,6078.75,0,35,19,19.53,4603,0,Somerset,1,1,Cable,38.606703,-120.58665900000001,1,94.55,2,6,Offer B,2958,1,0,1,0,65,0,1155.0,1269.45,0.0,6078.75,0,0,95684
1414,1,0,0,0,35,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,95.5,3418.2,0,27,59,45.62,3715,0,Sutter Creek,1,1,Fiber Optic,38.432145,-120.77068999999999,0,95.5,0,0,None,4610,1,0,0,0,35,1,2017.0,1596.6999999999996,0.0,3418.2,1,0,95685
1415,1,0,0,0,64,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),100.3,6603.8,0,51,2,9.95,4986,0,Thornton,0,1,Cable,38.157794,-121.520223,0,100.3,0,0,Offer B,1472,0,1,0,1,64,1,13.21,636.8,0.0,6603.8,0,1,95686
1416,0,0,1,1,58,0,No phone service,DSL,0,0,1,1,Two year,1,Credit card (automatic),55.5,3166.9,0,58,11,0.0,4080,0,Vacaville,1,0,Fiber Optic,38.333133000000004,-121.920151,1,55.5,0,1,Offer B,63157,1,0,1,1,58,1,348.0,0.0,0.0,3166.9,0,0,95687
1417,0,1,0,0,18,1,0,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),49.85,865.75,0,69,23,41.13,3283,0,Vacaville,0,0,Cable,38.419088,-122.02456799999999,0,49.85,0,0,None,32564,0,0,0,0,18,0,0.0,740.34,0.0,865.75,0,1,95688
1418,1,0,1,1,67,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),89.55,6373.1,0,38,53,6.15,6111,0,Volcano,0,1,Cable,38.481902000000005,-120.603668,1,89.55,3,4,Offer A,1273,0,0,1,1,67,0,3378.0,412.05,0.0,6373.1,0,0,95689
1419,1,0,1,1,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.15,1177.05,0,59,0,30.1,6373,0,Walnut Grove,0,1,NA,38.240419,-121.587535,1,19.15,3,2,None,2344,0,0,1,0,63,2,0.0,1896.3,0.0,1177.05,0,0,95690
1420,0,0,1,0,60,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.8,5985.75,0,22,51,34.48,6213,0,West Sacramento,0,0,DSL,38.627951,-121.59328700000002,1,99.8,0,9,None,19050,0,0,1,1,60,3,3053.0,2068.8,0.0,5985.75,1,0,95691
1421,1,1,0,0,9,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),84.4,732.5,1,67,20,30.8,5745,1,Wheatland,0,1,DSL,39.043387,-121.40983700000001,0,87.77600000000002,0,0,None,3600,0,0,0,0,9,8,146.0,277.2,0.0,732.5,0,0,95692
1422,0,0,1,1,70,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),113.05,7869.05,0,56,15,33.25,4203,0,Wilton,1,0,DSL,38.392559000000006,-121.22509299999999,1,113.05,2,4,Offer A,5889,1,0,1,1,70,0,1180.0,2327.5,0.0,7869.05,0,0,95693
1423,1,0,1,0,15,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.1,1504.05,1,62,32,40.7,2055,1,Winters,1,1,Cable,38.578604,-122.024579,1,105.144,0,1,None,8406,0,2,1,1,15,3,481.0,610.5,0.0,1504.05,0,0,95694
1424,0,0,0,1,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.95,936.7,0,32,0,9.19,3396,0,Woodland,0,0,NA,38.71967,-121.862416,0,19.95,0,0,None,38547,0,1,0,0,48,1,0.0,441.12,0.0,936.7,0,0,95695
1425,1,0,1,0,12,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,74.15,741.4,0,63,5,49.39,5426,0,Alta,1,1,Cable,39.218096,-120.79153000000001,1,74.15,0,7,None,751,1,0,1,1,12,1,37.0,592.6800000000002,0.0,741.4,0,0,95701
1426,1,1,1,0,71,1,1,Fiber optic,1,1,0,0,One year,1,Electronic check,92.0,6585.2,0,70,10,36.6,4322,0,Applegate,1,1,Fiber Optic,38.983388,-120.98881399999999,1,92.0,0,7,None,1526,1,0,1,0,71,0,65.85,2598.6,0.0,6585.2,0,1,95703
1427,1,1,0,0,44,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,73.85,3122.4,0,69,3,47.06,4374,0,Camino,1,1,Cable,38.748315999999996,-120.67551200000001,0,73.85,0,0,Offer B,4829,0,0,0,0,44,1,94.0,2070.640000000001,0.0,3122.4,0,0,95709
1428,1,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.45,50.45,1,37,10,28.25,2928,1,Colfax,0,1,DSL,39.084645,-120.89401399999998,0,52.468,0,0,None,8525,0,0,0,0,1,3,0.0,28.25,0.0,50.45,0,0,95713
1429,1,0,1,1,45,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.45,1088.25,0,43,0,47.31,3586,0,Dutch Flat,0,1,NA,39.197215,-120.83679,1,24.45,3,10,None,350,0,0,1,0,45,2,0.0,2128.9500000000007,0.0,1088.25,0,0,95714
1430,0,0,0,0,23,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),24.8,615.35,0,21,0,43.77,4402,0,Emigrant Gap,0,0,NA,39.23754,-120.720196,0,24.8,0,0,None,185,0,0,0,0,23,0,0.0,1006.71,0.0,615.35,1,0,95715
1431,0,0,1,0,43,1,1,DSL,0,0,1,0,One year,1,Bank transfer (automatic),64.85,2908.2,0,64,8,12.98,4000,0,Gold Run,0,0,Fiber Optic,39.170376,-120.838404,1,64.85,0,6,None,407,1,0,1,0,43,0,233.0,558.14,0.0,2908.2,0,0,95717
1432,1,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.75,739.9,0,49,0,17.92,5876,0,Kyburz,0,1,NA,38.766036,-120.209673,0,20.75,0,0,None,183,0,1,0,0,35,1,0.0,627.2,0.0,739.9,0,0,95720
1433,1,0,1,0,9,1,0,DSL,1,1,1,0,Month-to-month,1,Mailed check,68.95,593.85,0,47,7,34.64,2452,0,Echo Lake,0,1,Fiber Optic,38.851842,-120.076204,1,68.95,0,2,Offer E,69,1,0,1,0,9,2,0.0,311.76,0.0,593.85,0,1,95721
1434,1,0,0,0,12,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,99.95,1132.75,1,20,46,28.16,5598,1,Meadow Vista,0,1,Fiber Optic,39.003358,-121.022539,0,103.948,0,0,None,3747,1,3,0,1,12,5,0.0,337.92,0.0,1132.75,1,1,95722
1435,0,1,1,0,65,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),109.4,7227.45,0,68,29,15.3,4452,0,Pollock Pines,1,0,Fiber Optic,38.733908,-120.45341599999999,1,109.4,0,8,Offer B,8577,0,0,1,0,65,0,0.0,994.5,0.0,7227.45,0,1,95726
1436,0,0,0,0,2,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,91.4,193.6,1,50,8,39.62,5100,1,Soda Springs,1,0,Fiber Optic,39.279068,-120.414275,0,95.056,0,0,None,88,0,1,0,0,2,2,15.0,79.24,0.0,193.6,0,0,95728
1437,1,0,0,0,27,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,49.0,1291.35,0,61,15,2.69,5428,0,Twin Bridges,0,1,Cable,38.805481,-120.13287,0,49.0,0,0,None,25,0,2,0,0,27,1,194.0,72.63,0.0,1291.35,0,0,95735
1438,0,0,0,0,40,1,0,DSL,0,0,0,0,One year,1,Mailed check,50.25,2023.55,0,61,6,23.28,2449,0,Weimar,1,0,Fiber Optic,39.00978,-120.978273,0,50.25,0,0,None,31,0,0,0,0,40,0,121.0,931.2,0.0,2023.55,0,0,95736
1439,0,1,0,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.55,349.65,1,78,10,42.33,4028,1,Rancho Cordova,1,0,Cable,38.591134000000004,-121.161585,0,78.572,0,0,None,299,0,4,0,0,5,5,35.0,211.65,0.0,349.65,0,0,95742
1440,1,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.9,153.95,0,26,0,48.39,3152,0,Granite Bay,0,1,NA,38.749466,-121.184196,1,19.9,0,5,Offer E,20675,0,0,1,0,8,1,0.0,387.12,0.0,153.95,1,0,95746
1441,0,1,1,0,58,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),97.8,5458.8,0,66,28,45.37,6019,0,Roseville,0,0,Cable,38.784329,-121.373245,1,97.8,0,5,Offer B,25418,0,0,1,0,58,0,1528.0,2631.46,0.0,5458.8,0,0,95747
1442,0,0,1,1,52,1,0,Fiber optic,1,0,1,1,One year,0,Electronic check,100.3,5244.45,0,31,19,7.99,4811,0,Elk Grove,1,0,Fiber Optic,38.353629999999995,-121.44195,1,100.3,2,7,None,47065,0,0,1,1,52,0,996.0,415.48,0.0,5244.45,0,0,95758
1443,1,0,1,0,3,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,55.8,154.55,0,34,6,4.19,2662,0,El Dorado Hills,1,1,Fiber Optic,38.684437,-121.05563400000001,1,55.8,0,2,Offer E,22028,1,1,1,0,3,2,0.93,12.57,0.0,154.55,0,1,95762
1444,1,0,0,1,41,1,0,Fiber optic,1,1,1,1,Two year,1,Electronic check,111.15,4507.15,0,29,59,30.58,5038,0,Rocklin,1,1,Cable,38.823278,-121.281856,0,111.15,3,0,None,15494,1,0,0,1,41,2,2659.0,1253.78,0.0,4507.15,1,0,95765
1445,1,0,0,0,20,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,98.55,2031.95,0,26,59,23.22,3300,0,Woodland,0,1,DSL,38.694081,-121.69443100000001,0,98.55,0,0,None,15022,1,0,0,1,20,2,0.0,464.4,0.0,2031.95,1,1,95776
1446,1,0,0,1,1,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.05,50.05,0,24,69,43.05,5523,0,Sacramento,0,1,DSL,38.584505,-121.491956,0,50.05,3,0,Offer E,16599,0,0,0,0,1,1,0.0,43.05,0.0,50.05,1,1,95814
1447,1,0,0,1,4,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),80.8,332.45,1,28,84,42.33,5436,1,Sacramento,0,1,Fiber Optic,38.608405,-121.449942,0,84.03200000000001,0,0,None,25355,1,0,0,1,4,1,279.0,169.32,0.0,332.45,1,0,95815
1448,1,0,0,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.85,473.9,0,45,0,35.32,4263,0,Sacramento,0,1,NA,38.574856,-121.46503999999999,0,20.85,0,0,None,16164,0,0,0,0,23,0,0.0,812.36,0.0,473.9,0,0,95816
1449,0,1,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.5,106.8,0,67,0,2.03,3288,0,Sacramento,0,0,NA,38.550722,-121.457314,0,19.5,0,0,Offer E,14966,0,0,0,0,6,1,0.0,12.18,0.0,106.8,0,0,95817
1450,1,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.35,152.6,0,51,0,34.87,5416,0,Sacramento,0,1,NA,38.556306,-121.49581699999999,1,19.35,3,0,Offer E,21313,0,0,0,0,8,1,0.0,278.96,0.0,152.6,0,0,95818
1451,1,0,0,0,18,1,1,DSL,1,0,1,0,Month-to-month,0,Mailed check,69.5,1199.4,0,56,8,12.21,4466,0,Sacramento,1,1,DSL,38.567594,-121.43750700000001,0,69.5,0,0,None,15975,0,0,0,0,18,0,96.0,219.78000000000003,0.0,1199.4,0,0,95819
1452,1,1,0,0,52,0,No phone service,DSL,1,0,1,1,Month-to-month,1,Credit card (automatic),48.8,2555.05,0,69,19,0.0,4865,0,Sacramento,0,1,Fiber Optic,38.53508,-121.444144,0,48.8,0,0,Offer B,37031,0,0,0,1,52,2,0.0,0.0,0.0,2555.05,0,1,95820
1453,1,0,0,0,31,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,94.5,2979.2,0,56,18,45.92,3949,0,Sacramento,0,1,Fiber Optic,38.625096,-121.38365800000001,0,94.5,0,0,None,35426,0,0,0,1,31,1,53.63,1423.52,0.0,2979.2,0,1,95821
1454,1,0,1,1,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.65,654.85,0,20,0,24.64,4667,0,Sacramento,0,1,NA,38.512569,-121.49518400000001,1,20.65,1,5,None,44683,0,0,1,0,29,1,0.0,714.5600000000002,0.0,654.85,1,0,95822
1455,0,0,1,0,36,1,1,Fiber optic,1,1,0,1,Two year,1,Credit card (automatic),106.05,3834.4,0,54,18,19.24,4505,0,Sacramento,1,0,DSL,38.475465,-121.443625,1,106.05,0,4,None,72199,1,0,1,1,36,2,690.0,692.64,0.0,3834.4,0,0,95823
1456,0,0,1,0,16,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.0,1534.75,1,61,29,37.83,3794,1,Sacramento,0,0,Cable,38.517295000000004,-121.439819,1,104.0,0,1,None,30580,0,1,1,1,16,3,445.0,605.28,0.0,1534.75,0,0,95824
1457,1,0,1,0,42,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,108.3,4586.15,0,53,11,42.45,5106,0,Sacramento,1,1,Fiber Optic,38.590035,-121.41245500000001,1,108.3,0,1,None,30715,1,0,1,1,42,2,504.0,1782.9,0.0,4586.15,0,0,95825
1458,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.55,20.55,1,53,0,15.91,5636,1,Sacramento,0,1,NA,38.542532,-121.378826,0,20.55,0,0,None,38818,0,2,0,0,1,1,0.0,15.91,0.0,20.55,0,0,95826
1459,0,0,0,0,60,1,0,Fiber optic,0,1,1,1,Two year,1,Electronic check,99.65,5941.05,0,38,21,16.81,4616,0,Sacramento,1,0,Fiber Optic,38.549184999999994,-121.32838600000001,0,99.65,0,0,None,19611,0,0,0,1,60,0,1248.0,1008.6,0.0,5941.05,0,0,95827
1460,1,0,0,0,5,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,85.3,424.15,1,30,30,36.52,2264,1,Sacramento,1,1,Cable,38.486938,-121.39580500000001,0,88.712,0,0,None,54880,0,2,0,0,5,3,0.0,182.6,0.0,424.15,0,1,95828
1461,1,0,1,0,22,1,1,Fiber optic,1,0,1,0,Month-to-month,0,Credit card (automatic),95.9,2234.95,0,42,29,35.62,3207,0,Sacramento,0,1,Cable,38.486502,-121.334051,1,95.9,0,6,None,11396,1,0,1,0,22,0,0.0,783.64,0.0,2234.95,0,1,95829
1462,1,0,1,0,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.0,666.75,0,47,0,21.77,4175,0,Sacramento,0,1,NA,38.490508,-121.284171,1,20.0,0,7,None,592,0,0,1,0,36,1,0.0,783.72,0.0,666.75,0,0,95830
1463,0,0,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.4,281,1,19,46,41.12,4494,1,Sacramento,0,0,Fiber Optic,38.494832,-121.52944699999999,0,73.21600000000002,0,0,None,42832,0,3,0,1,4,4,129.0,164.48,0.0,281.0,1,0,95831
1464,1,0,0,0,9,1,0,DSL,1,0,0,1,Month-to-month,0,Mailed check,64.95,547.8,0,40,11,27.53,3013,0,Sacramento,0,1,Fiber Optic,38.445939,-121.49685500000001,0,64.95,0,0,Offer E,9063,1,0,0,1,9,3,0.0,247.77,0.0,547.8,0,1,95832
1465,1,0,1,1,1,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Credit card (automatic),74.6,74.6,0,28,59,42.99,5494,0,Sacramento,0,1,DSL,38.619049,-121.517552,1,74.6,1,5,None,31422,0,0,1,0,1,0,0.0,42.99,0.0,74.6,1,1,95833
1466,1,0,1,1,12,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.2,571.15,0,39,57,9.58,3582,0,Sacramento,0,1,Cable,38.646209000000006,-121.52446,1,49.2,3,8,Offer D,8403,0,0,1,0,12,0,0.0,114.96,0.0,571.15,0,1,95834
1467,0,0,0,0,23,1,1,DSL,0,0,1,1,One year,1,Mailed check,73.75,1756.6,0,37,3,35.03,3483,0,Sacramento,0,0,Cable,38.685069,-121.543709,0,73.75,0,0,Offer D,854,1,0,0,1,23,0,5.27,805.69,0.0,1756.6,0,1,95835
1468,1,0,0,0,62,1,1,Fiber optic,1,1,0,1,One year,1,Bank transfer (automatic),92.3,5731.45,0,35,16,24.35,6468,0,Sacramento,0,1,Cable,38.691607,-121.60228400000001,0,92.3,0,0,None,264,0,0,0,1,62,0,917.0,1509.7,0.0,5731.45,0,0,95837
1469,1,0,0,0,37,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),98.8,3475.55,1,27,46,30.72,3066,1,Sacramento,0,1,Fiber Optic,38.646096,-121.44243300000001,0,102.75200000000001,0,0,None,34894,1,0,0,1,37,0,1599.0,1136.64,0.0,3475.55,1,0,95838
1470,0,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.2,156.85,0,42,0,14.32,2879,0,Sacramento,0,0,NA,38.660441999999996,-121.346321,0,19.2,0,0,None,20993,0,0,0,0,8,2,0.0,114.56,0.0,156.85,0,0,95841
1471,1,0,1,0,31,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Credit card (automatic),88.65,2683.2,0,46,12,29.77,4821,0,Sacramento,1,1,Fiber Optic,38.687367,-121.34848000000001,1,88.65,0,9,None,31373,0,0,1,0,31,0,322.0,922.87,0.0,2683.2,0,0,95842
1472,1,0,1,1,13,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.4,896.75,1,36,23,2.92,3687,1,Antelope,0,1,Cable,38.715498,-121.36341100000001,1,77.376,0,1,None,36432,0,0,1,0,13,1,0.0,37.96,0.0,896.75,0,1,95843
1473,0,0,0,0,24,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.75,2407.3,1,35,20,37.69,4016,1,Sacramento,1,0,Cable,38.585826000000004,-121.376263,0,102.7,0,0,None,23362,0,1,0,1,24,2,481.0,904.56,0.0,2407.3,0,0,95864
1474,1,0,1,1,45,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),95.95,4456.65,0,54,19,22.31,5322,0,Marysville,1,1,Cable,39.19514,-121.503883,1,95.95,2,1,None,38091,0,0,1,1,45,0,0.0,1003.95,0.0,4456.65,0,1,95901
1475,0,1,1,0,69,1,1,Fiber optic,0,1,1,1,Two year,0,Credit card (automatic),105.4,6998.95,0,73,13,19.39,5467,0,Beale Afb,0,0,Cable,39.125310999999996,-121.392283,1,105.4,0,2,None,5654,1,0,1,1,69,0,0.0,1337.91,0.0,6998.95,0,1,95903
1476,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,36.8,0,35,0,15.83,5736,0,Alleghany,0,1,NA,39.467828000000004,-120.84138600000001,0,20.25,0,0,None,118,0,0,0,0,2,0,0.0,31.66,0.0,36.8,0,0,95910
1477,1,0,1,1,61,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,106.0,6547.7,1,52,23,46.95,4334,1,Arbuckle,0,1,Cable,38.982372999999995,-122.047751,1,110.24,0,1,None,4796,0,0,1,1,61,2,1506.0,2863.9500000000007,0.0,6547.7,0,0,95912
1478,1,0,0,0,41,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.7,4346.4,1,21,53,47.74,3316,1,Bangor,1,1,Cable,39.396584999999995,-121.38028999999999,0,108.88799999999999,0,0,None,626,0,1,0,1,41,4,2304.0,1957.34,0.0,4346.4,1,0,95914
1479,0,0,0,0,44,0,No phone service,DSL,0,0,1,1,One year,1,Electronic check,49.05,2265,0,58,3,0.0,3910,0,Berry Creek,1,0,Fiber Optic,39.657228,-121.37778,0,49.05,0,0,None,1279,0,0,0,1,44,2,0.0,0.0,0.0,2265.0,0,1,95916
1480,1,0,0,0,39,0,No phone service,DSL,0,0,0,0,One year,0,Mailed check,35.55,1309.15,0,41,14,0.0,3752,0,Biggs,1,1,Fiber Optic,39.457388,-121.818201,0,35.55,0,0,None,3169,1,0,0,0,39,0,183.0,0.0,0.0,1309.15,0,0,95917
1481,1,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,1,Credit card (automatic),65.1,4754.3,0,53,15,0.0,4969,0,Browns Valley,1,1,Fiber Optic,39.292334000000004,-121.32059699999999,1,65.1,0,7,Offer A,1477,1,1,1,1,72,3,713.0,0.0,0.0,4754.3,0,0,95918
1482,0,1,0,0,13,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.85,1235.55,0,74,24,26.68,3098,0,Brownsville,1,0,DSL,39.440687,-121.26358300000001,0,96.85,0,0,None,1237,0,0,0,1,13,0,0.0,346.84,0.0,1235.55,0,1,95919
1483,0,0,1,1,51,1,0,DSL,1,1,0,1,One year,1,Credit card (automatic),69.75,3562.5,0,50,14,17.95,5628,0,Butte City,0,0,Fiber Optic,39.449794,-121.93637199999999,1,69.75,0,2,None,303,1,0,1,1,51,0,0.0,915.45,0.0,3562.5,0,1,95920
1484,0,1,1,0,71,1,0,Fiber optic,0,1,1,1,Two year,1,Electronic check,99.2,7213.75,0,70,27,22.0,4951,0,Camptonville,1,0,Fiber Optic,39.432127,-121.09928700000002,1,99.2,0,6,None,632,0,1,1,1,71,2,0.0,1562.0,0.0,7213.75,0,1,95922
1485,1,1,0,0,22,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.7,2082.95,1,65,9,40.18,4458,1,Canyon Dam,0,1,Cable,40.171312,-121.120605,0,100.568,0,0,Offer D,86,0,0,0,1,22,1,187.0,883.96,0.0,2082.95,0,0,95923
1486,0,0,0,0,2,1,0,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),55.05,102.75,1,47,33,42.55,5855,1,Challenge,0,0,Fiber Optic,39.461768,-121.195825,0,57.251999999999995,0,0,Offer E,262,1,2,0,0,2,4,34.0,85.1,0.0,102.75,0,0,95925
1487,0,0,0,0,56,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,106.8,5914.4,0,49,2,32.43,6161,0,Chico,1,0,Fiber Optic,39.745712,-121.84333000000001,0,106.8,0,0,None,35808,0,0,0,1,56,0,118.0,1816.08,0.0,5914.4,0,0,95926
1488,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,51.25,51.25,0,32,26,39.3,4483,0,Chico,0,1,Fiber Optic,39.681488,-121.83721000000001,0,51.25,0,0,None,32848,0,0,0,0,1,3,0.0,39.3,0.0,51.25,0,1,95928
1489,0,0,1,1,23,1,0,DSL,1,1,0,0,One year,1,Mailed check,57.75,1282.85,0,30,41,12.88,3794,0,Clipper Mills,0,0,Fiber Optic,39.562239,-121.14836000000001,1,57.75,0,5,Offer D,282,1,0,1,0,23,0,0.0,296.24,0.0,1282.85,0,1,95930
1490,0,1,1,0,66,1,1,DSL,0,1,1,0,One year,1,Bank transfer (automatic),70.85,4738.85,0,73,17,44.01,5572,0,Colusa,1,0,Fiber Optic,39.273096,-122.05076299999999,1,70.85,0,0,None,7503,0,0,0,0,66,2,0.0,2904.66,0.0,4738.85,0,1,95932
1491,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.55,19.55,0,21,0,5.1,5750,0,Crescent Mills,0,0,NA,40.080342,-120.95780500000001,0,19.55,0,0,None,178,0,0,0,0,1,1,0.0,5.1,0.0,19.55,1,0,95934
1492,1,1,0,0,19,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,88.2,1775.8,1,74,10,39.97,5683,1,Dobbins,0,1,Cable,39.381174,-121.21191,0,91.728,0,0,Offer D,614,0,2,0,0,19,2,178.0,759.43,0.0,1775.8,0,0,95935
1493,1,0,0,0,11,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),79.5,795.65,0,20,52,8.48,2278,0,Downieville,1,1,Cable,39.578792,-120.780786,0,79.5,0,0,Offer D,404,0,0,0,0,11,0,414.0,93.28,0.0,795.65,1,0,95936
1494,0,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.75,145,1,44,0,46.13,2247,1,Dunnigan,0,0,NA,38.931425,-121.946081,1,19.75,0,1,Offer E,19,0,1,1,0,8,2,0.0,369.04,0.0,145.0,0,0,95937
1495,0,0,1,1,52,1,1,Fiber optic,1,1,0,1,Month-to-month,0,Bank transfer (automatic),98.15,4993.4,0,41,28,31.09,5123,0,Durham,1,0,Cable,39.607831,-121.77795900000001,1,98.15,1,6,None,3524,0,0,1,1,52,0,0.0,1616.68,0.0,4993.4,0,1,95938
1496,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.25,61.45,0,19,0,1.57,4050,0,Elk Creek,0,1,NA,39.53222,-122.594879,0,20.25,0,0,None,587,0,0,0,0,3,1,0.0,4.71,0.0,61.45,1,0,95939
1497,0,0,1,1,51,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Bank transfer (automatic),79.15,4018.55,0,29,71,2.53,6321,0,Forbestown,0,0,Fiber Optic,39.531028000000006,-121.24807,1,79.15,2,6,None,452,0,0,1,0,51,2,0.0,129.03,0.0,4018.55,1,1,95941
1498,1,1,0,0,15,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.65,1146.65,1,70,21,46.38,2099,1,Forest Ranch,0,1,DSL,40.077028000000006,-121.49416799999999,0,78.676,0,0,Offer D,1351,0,1,0,0,15,1,0.0,695.7,0.0,1146.65,0,1,95942
1499,1,1,1,0,64,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,94.25,6081.4,0,79,29,23.33,6020,0,Glenn,1,1,Fiber Optic,39.597975,-122.032248,1,94.25,0,9,Offer B,1454,0,0,1,0,64,0,0.0,1493.12,0.0,6081.4,0,1,95943
1500,0,0,0,0,37,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Credit card (automatic),40.2,1478.85,0,64,6,0.0,5924,0,Goodyears Bar,1,0,Fiber Optic,39.564113,-120.86883600000002,0,40.2,0,0,Offer C,76,0,1,0,1,37,1,89.0,0.0,0.0,1478.85,0,0,95944
1501,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.95,243.65,0,59,0,18.73,2884,0,Grass Valley,0,1,NA,39.194539,-120.98806599999999,0,19.95,0,0,Offer D,23990,0,0,0,0,13,0,0.0,243.49,0.0,243.65,0,0,95945
1502,1,0,1,0,49,1,1,DSL,1,0,0,0,One year,1,Electronic check,55.35,2633.95,0,29,52,42.19,5601,0,Penn Valley,0,1,Cable,39.203817,-121.19583999999999,1,55.35,0,3,None,9752,0,0,1,0,49,0,0.0,2067.31,0.0,2633.95,1,1,95946
1503,0,1,0,0,45,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),102.15,4735.35,0,74,15,34.12,5391,0,Greenville,1,0,Fiber Optic,40.160385999999995,-120.83542800000001,0,102.15,0,0,Offer B,2064,0,2,0,0,45,1,0.0,1535.4,0.0,4735.35,0,1,95947
1504,0,0,0,0,18,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.1,1247.75,0,19,26,2.76,4911,0,Gridley,0,0,Fiber Optic,39.346897999999996,-121.75953700000001,0,71.1,0,0,Offer D,9763,0,0,0,0,18,2,0.0,49.67999999999999,0.0,1247.75,1,1,95948
1505,1,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.7,74.7,1,69,22,11.34,3348,1,Grass Valley,0,1,DSL,39.099204,-121.13796200000002,0,77.688,0,0,None,17922,0,4,0,0,1,3,0.0,11.34,0.0,74.7,0,1,95949
1506,1,0,1,0,68,0,No phone service,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),54.1,3794.5,0,42,16,0.0,4601,0,Grimes,1,1,DSL,39.033058000000004,-121.89571799999999,1,54.1,0,7,Offer A,531,0,0,1,1,68,2,607.0,0.0,0.0,3794.5,0,0,95950
1507,1,0,0,0,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.65,1008.7,0,27,0,25.72,5708,0,Hamilton City,0,1,NA,39.732766999999996,-122.042298,0,19.65,0,0,None,1931,0,0,0,0,54,0,0.0,1388.88,0.0,1008.7,1,0,95951
1508,0,1,1,1,23,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),88.45,2130.55,0,74,53,2.03,3937,0,Live Oak,1,0,Fiber Optic,39.258746,-121.77696999999999,1,88.45,3,4,None,8695,0,0,1,0,23,1,0.0,46.69,0.0,2130.55,0,1,95953
1509,1,0,0,0,17,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.65,1313.55,1,62,8,30.61,3182,1,Magalia,1,1,Cable,39.933852,-121.58437099999999,0,79.71600000000002,0,0,None,11168,0,0,0,0,17,1,105.0,520.37,0.0,1313.55,0,0,95954
1510,1,0,1,0,71,1,1,DSL,1,1,0,1,Two year,0,Credit card (automatic),80.4,5727.15,0,22,41,18.04,5228,0,Maxwell,1,1,DSL,39.281194,-122.226568,1,80.4,0,2,Offer A,1146,1,0,1,1,71,0,2348.0,1280.84,0.0,5727.15,1,0,95955
1511,0,0,1,1,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.25,1372.9,0,56,0,48.75,5154,0,Meadow Valley,0,0,NA,39.937017,-121.058043,1,19.25,1,2,Offer A,301,0,0,1,0,67,2,0.0,3266.25,0.0,1372.9,0,0,95956
1512,0,0,1,1,14,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.8,1203.9,0,46,53,26.58,2452,0,Meridian,0,0,Cable,39.068071,-121.83263799999999,1,84.8,3,1,Offer D,776,0,0,1,0,14,0,638.0,372.12,0.0,1203.9,0,0,95957
1513,0,1,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,25.8,25.8,1,76,29,0.0,3884,1,Nevada City,0,0,DSL,39.333737,-120.858667,0,26.831999999999997,0,0,None,17269,0,1,0,0,1,2,0.0,0.0,0.0,25.8,0,1,95959
1514,0,0,0,1,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.5,1215.1,0,48,0,24.32,4370,0,North San Juan,0,0,NA,39.423046,-120.984472,0,19.5,1,0,None,565,0,0,0,0,63,1,0.0,1532.16,0.0,1215.1,0,0,95960
1515,0,0,0,0,41,1,1,DSL,0,0,0,1,One year,1,Electronic check,68.6,2877.05,0,36,30,36.93,4572,0,Olivehurst,1,0,Fiber Optic,39.082568,-121.55325,0,68.6,0,0,None,6439,1,0,0,1,41,1,0.0,1514.13,0.0,2877.05,0,1,95961
1516,0,0,1,0,17,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,92.6,1579.7,0,46,13,9.22,4756,0,Oregon House,0,0,DSL,39.342587,-121.24983300000001,1,92.6,0,10,Offer D,1519,0,0,1,1,17,1,0.0,156.74,0.0,1579.7,0,1,95962
1517,1,0,1,0,56,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,100.55,5514.95,0,28,48,46.9,4847,0,Orland,0,1,Fiber Optic,39.748037,-122.30216899999999,1,100.55,0,7,None,13706,0,0,1,1,56,0,2647.0,2626.4,0.0,5514.95,1,0,95963
1518,0,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.55,96.1,0,49,0,24.53,5967,0,Oroville,0,0,NA,39.624561,-121.552866,0,20.55,0,0,None,17782,0,0,0,0,5,1,0.0,122.65,0.0,96.1,0,0,95965
1519,0,0,0,0,2,0,No phone service,DSL,1,1,0,1,Month-to-month,1,Electronic check,42.6,72.4,1,49,23,0.0,4648,1,Oroville,0,0,DSL,39.473896,-121.415927,0,44.303999999999995,0,0,Offer E,28382,0,2,0,1,2,2,17.0,0.0,0.0,72.4,0,0,95966
1520,0,0,1,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.6,55.25,0,28,0,41.9,2941,0,Palermo,0,0,NA,39.435756,-121.552071,1,19.6,0,5,None,1254,0,0,1,0,3,0,0.0,125.7,0.0,55.25,1,0,95968
1521,1,0,0,0,37,1,1,DSL,1,1,0,0,One year,0,Electronic check,67.45,2443.3,0,42,14,13.04,5042,0,Paradise,1,1,DSL,39.69676,-121.644379,0,67.45,0,0,Offer C,28318,1,1,0,0,37,2,0.0,482.48,0.0,2443.3,0,1,95969
1522,0,0,0,0,29,1,0,DSL,1,1,0,1,Month-to-month,1,Bank transfer (automatic),68.85,1970.5,1,45,21,1.02,5449,1,Princeton,1,0,Cable,39.424957,-122.03930700000001,0,71.604,0,0,None,495,0,0,0,1,29,0,414.0,29.58,0.0,1970.5,0,0,95970
1523,1,0,0,0,8,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,43.55,335.4,0,44,23,7.02,3266,0,Quincy,0,1,Fiber Optic,39.971228,-121.04116599999999,0,43.55,0,0,None,6189,0,0,0,0,8,0,0.0,56.16,0.0,335.4,0,1,95971
1524,0,0,0,0,63,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),109.85,7002.95,0,40,20,19.01,5775,0,Chico,1,0,DSL,39.903271999999994,-121.843567,0,109.85,0,0,Offer B,26971,1,1,0,1,63,1,1401.0,1197.63,0.0,7002.95,0,0,95973
1525,0,0,1,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.65,158.95,0,61,0,5.01,4058,0,Richvale,0,0,NA,39.495768,-121.747472,1,20.65,1,7,None,74,0,0,1,0,7,4,0.0,35.07,0.0,158.95,0,0,95974
1526,0,0,0,0,3,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,95.4,293.15,0,52,28,17.01,2813,0,Rough And Ready,0,0,Fiber Optic,39.225634,-121.15616299999999,0,95.4,0,0,None,1601,0,1,0,1,3,1,82.0,51.03,0.0,293.15,0,0,95975
1527,1,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),21.0,1493.75,0,19,0,5.7,4974,0,Smartville,0,1,NA,39.176595,-121.291692,1,21.0,1,3,Offer A,963,0,0,1,0,72,1,0.0,410.4,0.0,1493.75,1,0,95977
1528,0,0,0,0,19,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,56.2,1093.4,0,57,22,40.22,3384,0,Stirling City,0,0,Cable,39.904002,-121.527823,0,56.2,0,0,Offer D,28,0,0,0,1,19,1,24.05,764.18,0.0,1093.4,0,1,95978
1529,0,0,1,0,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),18.4,1057.85,0,60,0,26.99,4375,0,Stonyford,0,0,NA,39.288127,-122.41584099999999,1,18.4,0,9,Offer B,844,0,0,1,0,59,0,0.0,1592.41,0.0,1057.85,0,0,95979
1530,1,0,1,1,2,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Credit card (automatic),90.0,190.05,1,51,8,46.92,3902,1,Strawberry Valley,1,1,Cable,39.584579999999995,-121.09325600000001,1,93.6,0,1,None,101,1,0,1,1,2,1,15.0,93.84,0.0,190.05,0,0,95981
1531,0,0,1,1,35,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,25.75,882.55,0,62,0,24.76,4194,0,Sutter,0,0,NA,39.172777,-121.80584499999999,1,25.75,1,5,Offer C,3193,0,2,1,0,35,1,0.0,866.6,0.0,882.55,0,0,95982
1532,1,0,0,0,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.6,300.4,0,64,0,8.54,2847,0,Taylorsville,0,1,NA,40.053684000000004,-120.74311599999999,0,19.6,0,0,Offer D,513,0,0,0,0,14,0,0.0,119.56,0.0,300.4,0,0,95983
1533,0,0,0,0,14,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.35,1025.95,1,42,22,18.74,4995,1,Twain,1,0,DSL,40.022184,-121.06238400000001,0,78.36399999999998,0,0,Offer D,73,0,0,0,0,14,0,226.0,262.36,0.0,1025.95,0,0,95984
1534,0,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.8,1436.95,0,29,0,8.39,5423,0,Washington,0,0,NA,39.34128,-120.78686699999999,1,19.8,2,7,Offer A,145,0,0,1,0,69,1,0.0,578.9100000000002,0.0,1436.95,1,0,95986
1535,1,1,1,0,7,1,1,DSL,1,1,0,0,Month-to-month,0,Electronic check,64.2,475,0,68,26,3.19,5116,0,Williams,0,1,Fiber Optic,39.117537,-122.284654,1,64.2,0,2,None,4579,1,0,1,0,7,0,12.35,22.33,0.0,475.0,0,1,95987
1536,1,0,1,1,69,1,0,DSL,1,1,1,0,Two year,1,Bank transfer (automatic),75.75,5388.15,0,64,18,44.33,5839,0,Willows,1,1,Fiber Optic,39.493990999999994,-122.286363,1,75.75,0,4,Offer A,8812,1,0,1,0,69,0,0.0,3058.77,0.0,5388.15,0,1,95988
1537,0,0,1,1,72,1,1,DSL,0,1,1,1,Two year,1,Electronic check,78.95,5730.15,0,56,6,26.04,5050,0,Yuba City,0,0,Fiber Optic,39.027409999999996,-121.61498200000001,1,78.95,0,10,Offer A,34967,1,0,1,1,72,0,0.0,1874.88,0.0,5730.15,0,1,95991
1538,1,0,0,0,8,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,100.85,819.55,1,56,7,3.27,3849,1,Yuba City,0,1,DSL,39.075694,-121.70606000000001,0,104.884,0,0,Offer E,27786,0,1,0,1,8,1,57.0,26.16,0.0,819.55,0,0,95993
1539,0,0,1,1,4,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,50.3,217.1,0,61,21,44.64,3147,0,Redding,0,0,Fiber Optic,40.587919,-122.46473200000001,1,50.3,1,8,None,31586,0,0,1,0,4,3,0.0,178.56,0.0,217.1,0,1,96001
1540,1,0,1,1,63,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),80.3,4896.35,0,30,48,18.88,5157,0,Redding,1,1,DSL,40.527834000000006,-122.318749,1,80.3,2,9,Offer B,30338,0,0,1,0,63,0,0.0,1189.4399999999996,0.0,4896.35,0,1,96002
1541,1,0,0,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.85,1434.1,0,52,0,3.43,4790,0,Redding,0,1,NA,40.677649,-122.29467,0,19.85,0,0,Offer A,41476,0,0,0,0,72,0,0.0,246.96,0.0,1434.1,0,0,96003
1542,0,0,0,0,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Electronic check,21.1,937.1,0,42,0,32.78,4791,0,Adin,0,0,NA,41.171578000000004,-120.91316100000002,0,21.1,0,0,Offer B,615,0,0,0,0,46,1,0.0,1507.88,0.0,937.1,0,0,96006
1543,0,0,1,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.95,330.15,1,55,11,17.08,2969,1,Anderson,0,0,Cable,40.448632,-122.306657,1,72.748,0,1,Offer E,21418,0,1,1,0,5,1,0.0,85.39999999999998,0.0,330.15,0,1,96007
1544,1,0,1,0,30,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.0,1474.9,0,53,6,23.16,4715,0,Bella Vista,1,1,Cable,40.722733000000005,-122.10966599999999,1,50.0,0,10,Offer C,899,0,0,1,0,30,1,88.0,694.8,0.0,1474.9,0,0,96008
1545,1,0,0,0,63,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),104.75,6536.5,0,52,21,48.75,5882,0,Bieber,1,1,Cable,41.083464,-121.107929,0,104.75,0,0,Offer B,595,0,1,0,1,63,1,0.0,3071.25,0.0,6536.5,0,1,96009
1546,0,0,0,0,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.85,1128.1,0,53,0,31.12,6213,0,Big Bar,0,0,NA,40.775271999999994,-123.28741399999998,0,19.85,0,0,Offer B,269,0,0,0,0,60,0,0.0,1867.2,0.0,1128.1,0,0,96010
1547,0,0,1,0,63,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,107.5,6873.75,1,50,23,1.93,6144,1,Big Bend,1,0,DSL,41.096569,-121.87908200000001,1,111.8,0,1,None,265,0,0,1,1,63,3,1581.0,121.59,0.0,6873.75,0,0,96011
1548,1,0,1,1,25,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,85.9,2199.05,0,26,59,11.79,3153,0,Burney,0,1,Cable,40.946785,-121.719489,1,85.9,3,0,Offer C,4552,1,0,0,0,25,4,0.0,294.75,0.0,2199.05,1,1,96013
1549,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.85,45.85,1,58,13,44.75,5930,1,Callahan,0,1,Cable,41.388397,-122.79463600000001,0,47.68400000000001,0,0,Offer E,290,0,0,0,0,1,3,0.0,44.75,0.0,45.85,0,0,96014
1550,1,1,1,0,6,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,80.8,457.1,0,75,17,16.87,5611,0,Canby,1,1,Fiber Optic,41.486953,-120.913975,1,80.8,0,4,None,417,0,0,1,0,6,0,0.0,101.22,0.0,457.1,0,1,96015
1551,1,0,0,0,22,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.25,566.5,0,61,0,4.79,3403,0,Cassel,0,1,NA,40.936285,-121.57269199999999,0,25.25,0,0,Offer D,344,0,0,0,0,22,0,0.0,105.38,0.0,566.5,0,0,96016
1552,0,0,1,1,31,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),80.55,2471.6,0,58,2,28.52,3491,0,Castella,0,0,Fiber Optic,41.121108,-122.33661299999999,1,80.55,0,9,Offer C,228,1,0,1,1,31,1,49.0,884.12,0.0,2471.6,0,0,96017
1553,0,0,1,1,39,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),81.5,3107.3,0,64,76,40.68,2042,0,Shasta Lake,1,0,DSL,40.692523,-122.369876,1,81.5,5,7,Offer C,6277,1,0,1,0,39,0,0.0,1586.52,0.0,3107.3,0,1,96019
1554,1,0,0,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.9,518.3,0,31,0,31.73,5895,0,Chester,0,1,NA,40.243494,-121.15473300000001,0,20.9,0,0,Offer C,2664,0,0,0,0,26,0,0.0,824.98,0.0,518.3,0,0,96020
1555,0,0,1,0,53,1,0,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),106.1,5769.75,1,44,12,30.09,4471,1,Corning,1,0,DSL,39.913777,-122.289984,1,110.344,0,1,None,13840,0,0,1,1,53,3,692.0,1594.77,0.0,5769.75,0,0,96021
1556,0,0,0,0,1,1,0,Fiber optic,0,1,1,0,Month-to-month,0,Electronic check,91.7,91.7,1,20,57,17.23,4319,1,Cottonwood,0,0,Cable,40.336392,-122.44853300000001,0,95.368,0,0,Offer E,12348,1,0,0,1,1,3,0.0,17.23,0.0,91.7,1,1,96022
1557,1,0,0,0,12,1,1,DSL,1,1,0,0,Month-to-month,1,Electronic check,67.25,832.3,0,54,4,45.8,4334,0,Dorris,0,1,Cable,41.949216,-122.05006200000001,0,67.25,0,0,Offer D,1162,1,0,0,0,12,1,3.33,549.5999999999998,0.0,832.3,0,1,96023
1558,0,0,0,0,16,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),95.6,1555.65,1,39,33,18.99,5915,1,Douglas City,1,0,Cable,40.586588,-122.903677,0,99.424,0,0,Offer D,960,0,0,0,1,16,1,513.0,303.84,0.0,1555.65,0,0,96024
1559,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,45.3,0,52,0,25.92,5994,0,Dunsmuir,0,0,NA,41.212695000000004,-122.392067,0,20.35,0,0,None,2602,0,0,0,0,2,3,0.0,51.84,0.0,45.3,0,0,96025
1560,1,0,0,1,39,0,No phone service,DSL,1,0,1,0,One year,0,Bank transfer (automatic),45.05,1790.6,0,40,13,0.0,4003,0,Etna,0,1,Fiber Optic,41.405193,-123.008567,0,45.05,0,0,Offer C,2156,1,0,0,0,39,0,0.0,0.0,0.0,1790.6,0,1,96027
1561,1,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.95,74.95,1,59,29,30.07,2591,1,Fall River Mills,0,1,Cable,41.017282,-121.46894499999999,0,77.94800000000002,0,0,Offer E,1902,0,4,0,0,1,2,0.0,30.07,0.0,74.95,0,0,96028
1562,0,0,1,1,7,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,34.65,246.6,0,37,17,0.0,5996,0,Flournoy,0,0,DSL,39.847840000000005,-122.544556,1,34.65,1,8,None,84,1,0,1,0,7,1,42.0,0.0,0.0,246.6,0,0,96029
1563,1,1,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.35,261.65,0,77,25,30.11,4140,0,Forks Of Salmon,0,1,Fiber Optic,41.232128,-123.194748,0,69.35,0,0,None,170,0,0,0,0,4,0,6.54,120.44,0.0,261.65,0,1,96031
1564,1,1,0,0,10,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.35,898.35,1,71,15,41.37,5353,1,Escondido,0,1,Cable,33.141265000000004,-116.967221,0,99.164,0,0,Offer D,48690,0,0,0,0,10,1,135.0,413.7,0.0,898.35,0,0,92027
1565,0,0,0,0,55,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,81.55,4509.5,0,39,4,22.34,5167,0,French Gulch,1,0,Fiber Optic,40.740138,-122.587476,0,81.55,0,0,Offer B,373,0,0,0,0,55,0,0.0,1228.7,0.0,4509.5,0,1,96033
1566,1,0,1,1,72,1,0,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),75.4,5480.25,0,43,18,42.16,4171,0,Gazelle,1,1,Fiber Optic,41.411315,-122.697236,1,75.4,0,7,None,392,0,0,1,1,72,0,0.0,3035.5199999999995,0.0,5480.25,0,1,96034
1567,0,0,1,0,10,1,0,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),67.8,653.15,0,62,7,37.08,2709,0,Gerber,1,0,Cable,40.031940000000006,-122.176023,1,67.8,0,6,Offer D,3357,0,0,1,1,10,1,0.0,370.8,0.0,653.15,0,1,96035
1568,1,1,0,0,11,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,111.4,1183.05,0,75,13,2.63,3175,0,Greenview,1,1,Fiber Optic,41.528541,-122.955018,0,111.4,0,0,None,295,1,2,0,0,11,2,154.0,28.93,0.0,1183.05,0,0,96037
1569,0,0,1,1,15,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,46.3,639.45,0,24,27,24.27,3103,0,Grenada,0,0,DSL,41.599978,-122.539381,1,46.3,3,7,Offer D,616,0,0,1,0,15,0,173.0,364.05,0.0,639.45,1,0,96038
1570,0,0,1,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.4,478.75,0,48,0,39.59,4698,0,Happy Camp,0,0,NA,41.831901,-123.487478,1,20.4,1,1,Offer D,1294,0,0,1,0,23,1,0.0,910.57,0.0,478.75,0,0,96039
1571,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,20.05,0,46,0,7.66,4221,0,Hat Creek,0,1,NA,40.789799,-121.474529,0,20.05,3,0,None,397,0,0,0,0,1,0,0.0,7.66,0.0,20.05,0,0,96040
1572,0,1,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.0,127.1,1,76,7,30.14,4145,1,Fallbrook,0,0,DSL,33.362575,-117.299644,0,46.8,0,0,None,42239,0,0,0,0,3,3,9.0,90.42,0.0,127.1,0,0,92028
1573,1,0,1,1,47,1,0,Fiber optic,1,1,0,1,One year,1,Electronic check,96.1,4391.45,0,23,52,15.59,5793,0,Hornbrook,1,1,DSL,41.962127,-122.52769599999999,1,96.1,2,1,Offer B,1026,0,2,1,1,47,1,228.36,732.73,0.0,4391.45,1,1,96044
1574,0,0,0,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.65,270.6,0,36,0,23.56,4818,0,Hyampom,0,0,NA,40.648024,-123.465088,0,19.65,0,0,None,268,0,0,0,0,15,0,0.0,353.4,0.0,270.6,0,0,96046
1575,1,0,0,0,66,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,99.5,6710.5,1,62,29,25.82,4001,1,Igo,1,1,Cable,40.524535,-122.647172,0,103.48,0,0,Offer A,911,0,0,0,1,66,4,194.6,1704.12,0.0,6710.5,0,1,96047
1576,0,1,1,0,68,1,0,DSL,0,1,0,0,One year,1,Bank transfer (automatic),60.65,3975.9,0,78,20,40.55,6418,0,Junction City,1,0,DSL,40.913191999999995,-123.06597,1,60.65,0,2,None,734,1,0,1,0,68,0,0.0,2757.4,0.0,3975.9,0,1,96048
1577,0,0,1,1,17,1,0,Fiber optic,0,0,1,1,One year,0,Bank transfer (automatic),98.6,1704.95,1,38,9,5.4,5160,1,Klamath River,1,0,DSL,41.816595,-122.94828700000001,1,102.544,0,1,Offer D,482,1,2,1,1,17,3,153.0,91.8,0.0,1704.95,0,0,96050
1578,0,0,0,0,7,1,0,DSL,0,0,1,0,Month-to-month,1,Mailed check,59.5,415.95,1,54,24,2.24,4661,1,Lakehead,0,0,Cable,40.883853,-122.41825800000001,0,61.88,0,0,Offer E,1236,1,0,0,0,7,6,100.0,15.68,0.0,415.95,0,0,96051
1579,1,1,1,0,12,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.45,950.2,1,77,21,6.97,5374,1,Lewiston,0,1,Cable,40.704293,-122.803899,1,83.66799999999999,0,1,Offer D,1845,0,0,1,0,12,1,200.0,83.64,0.0,950.2,0,0,96052
1580,0,1,1,0,21,1,1,DSL,0,1,0,1,One year,0,Bank transfer (automatic),71.7,1497.05,0,73,18,30.3,2784,0,Lookout,1,0,Fiber Optic,41.280478,-121.160249,1,71.7,0,4,None,386,0,0,1,0,21,0,0.0,636.3000000000002,0.0,1497.05,0,1,96054
1581,1,0,0,0,21,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Mailed check,36.0,780.15,0,39,9,0.0,3378,0,Los Molinos,0,1,DSL,40.059385,-122.091481,0,36.0,0,0,None,3756,1,0,0,0,21,0,70.0,0.0,0.0,780.15,0,0,96055
1582,0,0,1,1,56,1,1,DSL,1,0,1,0,One year,0,Bank transfer (automatic),65.2,3512.15,0,62,11,39.72,4775,0,Mcarthur,0,0,Cable,41.108309999999996,-121.36036200000001,1,65.2,0,1,Offer B,1554,0,0,1,0,56,3,386.0,2224.32,0.0,3512.15,0,0,96056
1583,0,0,1,1,6,1,1,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),48.95,273.25,0,28,82,24.83,3061,0,Mccloud,0,0,Fiber Optic,41.251321999999995,-122.105209,1,48.95,1,1,Offer E,1586,0,0,1,0,6,1,0.0,148.98,0.0,273.25,1,1,96057
1584,0,1,0,0,65,0,No phone service,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),53.5,3517.9,0,75,9,0.0,5693,0,Macdoel,1,0,Fiber Optic,41.769709000000006,-121.92063,0,53.5,0,0,Offer B,816,0,0,0,0,65,0,317.0,0.0,0.0,3517.9,0,0,96058
1585,1,0,1,0,42,1,1,DSL,1,0,1,1,One year,0,Credit card (automatic),80.45,3375.9,0,30,82,17.31,4397,0,Manton,0,1,Cable,40.426679,-121.850421,1,80.45,0,1,Offer B,598,1,0,1,1,42,0,2768.0,727.02,0.0,3375.9,0,0,96059
1586,0,0,1,1,68,1,1,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),109.05,7508.55,0,55,53,18.42,6391,0,Mill Creek,1,0,Cable,40.331975,-121.460674,1,109.05,3,1,None,78,1,0,1,1,68,0,3980.0,1252.5600000000004,0.0,7508.55,0,0,96061
1587,1,0,1,1,48,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),26.3,1245.05,0,59,0,20.73,2111,0,Millville,0,1,NA,40.531257000000004,-122.14813899999999,1,26.3,3,1,Offer B,830,0,0,1,0,48,2,0.0,995.04,0.0,1245.05,0,0,96062
1588,0,1,0,0,50,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,106.8,5347.95,0,66,14,10.6,5746,0,Mineral,0,0,Fiber Optic,40.408796,-121.579609,0,106.8,0,0,Offer B,124,1,0,0,0,50,0,74.87,530.0,0.0,5347.95,0,1,96063
1589,0,1,0,0,7,1,0,DSL,0,1,1,0,Month-to-month,1,Electronic check,64.95,493.65,0,67,7,7.82,4615,0,Fallbrook,1,0,Cable,33.362575,-117.299644,0,64.95,0,0,None,42239,0,0,0,0,7,0,35.0,54.74,0.0,493.65,0,0,92028
1590,0,0,1,1,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,19.35,1263.85,0,31,0,41.84,4566,0,Montgomery Creek,0,0,NA,40.877552,-121.885884,1,19.35,3,0,Offer B,431,0,0,0,0,63,1,0.0,2635.92,0.0,1263.85,0,0,96065
1591,1,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),21.1,385.55,0,24,0,34.02,2842,0,Mount Shasta,0,1,NA,41.33832,-122.290756,0,21.1,0,0,None,7309,0,0,0,0,17,0,0.0,578.34,0.0,385.55,1,0,96067
1592,0,0,1,1,42,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),77.95,3384,1,53,20,34.02,5396,1,Nubieber,0,0,Cable,41.082471999999996,-121.19521499999999,1,81.06800000000001,0,1,None,240,0,1,1,0,42,2,677.0,1428.84,0.0,3384.0,0,0,96068
1593,1,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,18.85,84.2,0,41,0,39.04,5279,0,Oak Run,0,1,NA,40.689243,-122.037023,1,18.85,1,1,Offer E,829,0,0,1,0,4,0,0.0,156.16,0.0,84.2,0,0,96069
1594,0,0,0,1,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),26.0,1638.7,0,51,0,2.83,4535,0,Old Station,0,0,NA,40.656287,-121.42896499999999,0,26.0,3,0,Offer B,182,0,0,0,0,62,0,0.0,175.46,0.0,1638.7,0,0,96071
1595,1,1,0,0,2,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.7,165.4,1,74,12,6.51,2803,1,Palo Cedro,0,1,DSL,40.582399,-122.19551200000001,0,77.688,0,0,None,4931,0,1,0,0,2,1,0.0,13.02,0.0,165.4,0,1,96073
1596,0,0,1,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.35,120.25,0,45,22,7.7,4917,0,Paskenta,0,0,Cable,39.884395,-122.58751299999999,1,70.35,0,1,Offer E,263,0,0,1,0,2,0,2.65,15.4,0.0,120.25,0,1,96074
1597,1,0,1,0,48,1,1,Fiber optic,1,1,1,0,Two year,1,Bank transfer (automatic),96.9,4473.45,0,33,18,6.1,2613,0,Paynes Creek,1,1,Cable,40.343213,-121.81541200000001,1,96.9,0,1,Offer B,433,0,2,1,0,48,2,0.0,292.7999999999999,0.0,4473.45,0,1,96075
1598,1,0,1,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.55,520.55,0,53,0,44.19,4430,0,Platina,0,1,NA,40.367964,-122.937379,1,19.55,0,1,Offer C,215,0,1,1,0,27,1,0.0,1193.13,0.0,520.55,0,0,96076
1599,0,0,1,1,70,1,0,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),80.4,5717.85,0,28,52,39.78,6367,0,Red Bluff,1,0,Fiber Optic,40.186772,-122.388361,1,80.4,0,4,None,26438,1,0,1,1,70,0,2973.0,2784.6,0.0,5717.85,1,0,96080
1600,1,1,0,0,1,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,88.8,88.8,1,77,22,49.6,3106,1,Round Mountain,1,1,Cable,40.923558,-122.059933,0,92.352,0,0,None,459,0,0,0,0,1,1,0.0,49.6,0.0,88.8,0,0,96084
1601,1,0,1,0,46,1,1,Fiber optic,0,1,1,0,One year,1,Electronic check,94.65,4312.5,0,44,3,10.13,4120,0,Scott Bar,1,1,Cable,41.737961999999996,-123.07557,1,94.65,0,1,Offer B,88,0,0,1,0,46,0,129.0,465.98,0.0,4312.5,0,0,96085
1602,1,0,0,0,30,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.25,2755.35,1,33,21,30.06,5654,1,San Diego,0,1,Cable,32.957195,-117.202542,0,93.86,0,0,None,28201,0,2,0,1,30,1,579.0,901.8,0.0,2755.35,0,0,92130
1603,0,0,0,0,15,1,1,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),64.65,994.55,1,51,29,47.57,4780,1,San Diego,0,0,DSL,32.957195,-117.202542,0,67.236,0,0,Offer D,28201,0,0,0,1,15,1,28.84,713.55,0.0,994.55,0,1,92130
1604,1,0,1,1,69,1,1,Fiber optic,0,1,1,0,One year,0,Credit card (automatic),95.75,6511.25,0,35,27,42.45,5561,0,Shingletown,1,1,Fiber Optic,40.497440999999995,-121.827524,1,95.75,2,9,None,4231,0,0,1,0,69,0,0.0,2929.05,0.0,6511.25,0,1,96088
1605,1,0,0,0,65,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.55,1218.65,0,34,0,44.7,4309,0,Tehama,0,1,NA,40.021786999999996,-122.127576,0,19.55,0,0,Offer B,405,0,0,0,0,65,0,0.0,2905.5,0.0,1218.65,0,0,96090
1606,1,1,1,1,72,1,0,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),104.1,7447.7,0,67,25,16.82,5092,0,Trinity Center,1,1,Fiber Optic,41.081846999999996,-122.70054499999999,1,104.1,2,4,None,734,1,0,1,0,72,0,0.0,1211.04,0.0,7447.7,0,1,96091
1607,1,1,1,0,13,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),89.05,1169.35,1,76,6,1.47,3861,1,San Diego,0,1,Cable,32.957195,-117.202542,1,92.61200000000001,0,1,Offer D,28201,1,0,1,0,13,1,70.0,19.11,0.0,1169.35,0,0,92130
1608,1,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.1,279.5,0,46,0,31.6,2185,0,Weaverville,0,1,NA,40.759401000000004,-122.93933700000001,0,20.1,0,0,None,3749,0,0,0,0,17,0,0.0,537.2,0.0,279.5,0,0,96093
1609,1,0,1,0,51,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,111.55,5720.35,0,23,76,39.32,4053,0,Weed,1,1,Fiber Optic,41.465121,-122.38094699999999,1,111.55,0,2,Offer B,5896,1,0,1,1,51,2,4347.0,2005.32,0.0,5720.35,1,0,96094
1610,1,0,1,1,51,1,0,DSL,1,1,0,0,Two year,0,Credit card (automatic),60.5,3121.45,0,40,10,9.53,4994,0,Whitmore,0,1,Cable,40.637105,-121.906949,1,60.5,0,5,Offer B,843,1,0,1,0,51,1,0.0,486.03,0.0,3121.45,0,1,96096
1611,0,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),90.95,6468.6,0,52,15,42.64,6091,0,Yreka,1,0,DSL,41.764869,-122.67131599999999,1,90.95,0,6,None,9538,1,0,1,1,72,1,97.03,3070.08,0.0,6468.6,0,1,96097
1612,1,0,1,1,67,1,1,Fiber optic,0,1,0,0,One year,0,Electronic check,87.4,5918.8,1,34,11,28.4,4421,1,San Diego,1,1,Fiber Optic,32.957195,-117.202542,1,90.89600000000002,0,1,Offer A,28201,0,0,1,0,67,0,651.0,1902.8,0.0,5918.8,0,0,92130
1613,1,0,0,0,34,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.7,675.6,0,31,0,36.52,4136,0,Blairsden Graeagle,0,1,NA,39.783747,-120.661032,0,19.7,0,0,Offer C,1839,0,0,0,0,34,1,0.0,1241.68,0.0,675.6,0,0,96103
1614,1,0,1,0,67,0,No phone service,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),50.95,3521.7,0,39,6,0.0,6395,0,Cedarville,0,1,Fiber Optic,41.505916,-120.152505,1,50.95,0,10,None,857,1,0,1,1,67,0,211.0,0.0,0.0,3521.7,0,0,96104
1615,0,0,1,0,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.05,923.1,0,56,0,22.1,5579,0,Chilcoot,0,0,NA,39.872961,-120.198876,1,20.05,0,3,None,650,0,0,1,0,49,1,0.0,1082.9,0.0,923.1,0,0,96105
1616,1,0,1,1,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.4,1110.35,0,38,0,25.32,4497,0,Clio,0,1,NA,39.745805,-120.580882,1,19.4,3,8,None,88,0,0,1,0,53,0,0.0,1341.96,0.0,1110.35,0,0,96106
1617,1,0,0,0,27,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,59.45,1611.65,0,55,25,33.94,4818,0,Coleville,1,1,Fiber Optic,38.42528,-119.47574099999999,0,59.45,0,0,None,1332,1,0,0,0,27,1,403.0,916.38,0.0,1611.65,0,0,96107
1618,0,1,0,0,23,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,94.75,2293.6,1,77,25,31.17,2740,1,San Diego,0,0,Fiber Optic,32.957195,-117.202542,0,98.54,0,0,Offer D,28201,0,1,0,0,23,4,573.0,716.9100000000002,0.0,2293.6,0,0,92130
1619,1,0,0,0,69,1,1,DSL,1,1,0,1,Two year,1,Credit card (automatic),81.5,5553.25,0,46,26,3.24,5286,0,Doyle,1,1,Fiber Optic,40.012675,-120.10185700000001,0,81.5,0,0,None,1177,1,0,0,1,69,0,0.0,223.56,0.0,5553.25,0,1,96109
1620,0,0,1,1,2,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),29.05,44.75,0,51,27,0.0,4998,0,Eagleville,0,0,Fiber Optic,41.280341,-120.15038100000001,1,29.05,2,4,Offer E,132,1,0,1,0,2,1,0.0,0.0,0.0,44.75,0,1,96110
1621,0,0,0,0,35,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.45,3029.1,1,32,19,19.07,5874,1,San Diego,0,0,DSL,32.957195,-117.202542,0,89.90799999999999,0,0,None,28201,0,2,0,0,35,3,576.0,667.45,0.0,3029.1,0,0,92130
1622,0,0,1,0,46,1,0,DSL,1,1,0,1,One year,0,Mailed check,70.6,3231.05,0,45,27,44.75,5433,0,Herlong,0,0,Fiber Optic,40.198234,-120.18088999999999,1,70.6,0,6,None,946,1,0,1,1,46,4,0.0,2058.5,0.0,3231.05,0,1,96113
1623,0,0,0,0,54,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),97.2,5129.45,0,39,8,31.55,4971,0,Janesville,0,0,DSL,40.294034,-120.512622,0,97.2,0,0,None,3093,0,0,0,1,54,2,0.0,1703.7,0.0,5129.45,0,1,96114
1624,0,0,1,0,56,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,98.25,5508.35,1,21,53,19.16,4886,1,San Diego,0,0,Cable,32.957195,-117.202542,1,102.18,0,1,None,28201,0,0,1,1,56,1,2919.0,1072.96,0.0,5508.35,1,0,92130
1625,0,0,1,0,9,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.75,655.9,1,46,28,31.75,5105,1,San Diego,1,0,Cable,32.957195,-117.202542,1,78.78,0,1,Offer E,28201,0,0,1,0,9,4,184.0,285.75,0.0,655.9,0,0,92130
1626,1,0,0,0,20,1,1,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),59.2,1191.2,0,53,17,33.14,5924,0,Litchfield,0,1,DSL,40.507272,-120.338228,0,59.2,0,0,None,385,1,0,0,0,20,0,0.0,662.8,0.0,1191.2,0,1,96117
1627,1,0,0,0,11,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,75.9,866.4,0,20,27,13.55,4278,0,Loyalton,0,1,Fiber Optic,39.637471000000005,-120.22633799999998,0,75.9,0,0,None,1822,0,0,0,0,11,3,0.0,149.05,0.0,866.4,1,1,96118
1628,0,1,1,0,30,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,90.05,2627.2,0,68,27,47.75,3792,0,Madeline,0,0,DSL,41.042003,-120.50608600000001,1,90.05,0,8,Offer C,85,0,0,1,0,30,0,0.0,1432.5,0.0,2627.2,0,1,96119
1629,1,0,1,0,68,1,0,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),70.95,4741.45,0,56,3,11.94,5036,0,Markleeville,1,1,DSL,38.735789000000004,-119.85798,1,70.95,0,4,None,957,0,0,1,1,68,2,142.0,811.92,0.0,4741.45,0,0,96120
1630,1,1,1,0,38,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,102.6,4009.2,0,79,24,4.75,5469,0,Milford,1,1,Fiber Optic,40.181278999999996,-120.392967,1,102.6,0,7,Offer C,481,0,0,1,0,38,3,962.0,180.5,45.81,4009.2,0,0,96121
1631,0,1,1,0,17,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),85.35,1463.45,1,80,7,36.82,3209,1,San Diego,1,0,Fiber Optic,32.957195,-117.202542,1,88.764,0,1,Offer D,28201,0,0,1,0,17,1,102.0,625.94,0.0,1463.45,0,0,92130
1632,1,0,0,0,48,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),106.1,5082.8,1,55,4,24.73,5898,1,San Diego,1,1,Cable,32.957195,-117.202542,0,110.344,0,0,None,28201,0,2,0,1,48,5,203.0,1187.04,0.0,5082.8,0,0,92130
1633,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,43.8,43.8,0,39,3,37.5,4633,0,Calpine,0,0,Fiber Optic,39.672813,-120.456699,0,43.8,0,0,Offer E,322,0,0,0,0,1,0,0.0,37.5,0.0,43.8,0,1,96124
1634,1,0,1,1,63,0,No phone service,DSL,1,1,1,1,Two year,0,Electronic check,59.0,3707.6,0,36,5,0.0,5639,0,Sierra City,1,1,Fiber Optic,39.600599,-120.636358,1,59.0,0,1,None,348,0,0,1,1,63,2,0.0,0.0,0.0,3707.6,0,1,96125
1635,0,0,0,0,3,1,0,DSL,0,0,1,1,One year,1,Electronic check,69.95,220.45,0,58,17,29.51,2754,0,Sierraville,1,0,DSL,39.559709000000005,-120.34563899999999,0,69.95,0,0,Offer E,227,0,0,0,1,3,0,37.0,88.53,0.0,220.45,0,0,96126
1636,0,0,0,0,48,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),24.35,1133.7,0,25,0,13.67,4200,0,Standish,0,0,NA,40.346634,-120.386422,0,24.35,0,0,None,408,0,0,0,0,48,2,0.0,656.16,0.0,1133.7,1,0,96128
1637,1,0,0,0,66,0,No phone service,DSL,0,0,0,0,One year,0,Credit card (automatic),29.45,1983.15,0,45,15,0.0,5112,0,Susanville,0,1,Fiber Optic,40.559177000000005,-120.612113,0,29.45,0,0,None,19440,1,0,0,0,66,0,0.0,0.0,0.0,1983.15,0,1,96130
1638,0,0,1,1,68,1,1,Fiber optic,0,1,0,0,Two year,1,Credit card (automatic),84.4,5746.75,0,44,30,24.94,5045,0,Termo,1,0,Fiber Optic,41.027281,-120.669427,1,84.4,1,3,None,72,0,0,1,0,68,0,1724.0,1695.92,0.0,5746.75,0,0,96132
1639,1,1,0,0,17,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.05,770.6,1,68,2,40.93,3797,1,San Diego,0,1,Fiber Optic,32.957195,-117.202542,0,46.852,0,0,None,28201,0,0,0,0,17,0,0.0,695.81,0.0,770.6,0,1,92130
1640,0,0,1,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.65,134.05,0,20,0,41.64,3575,0,Tulelake,0,0,NA,41.813521,-121.49266599999999,1,20.65,0,2,Offer E,2595,0,0,1,0,7,0,0.0,291.48,0.0,134.05,1,0,96134
1641,1,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),87.1,6230.1,0,48,26,12.02,5993,0,Wendel,1,1,Cable,40.345949,-120.08118700000001,1,87.1,0,5,None,162,1,0,1,1,72,0,0.0,865.4399999999998,0.0,6230.1,0,1,96136
1642,0,0,1,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,573.05,0,46,0,5.69,2712,0,Westwood,0,0,NA,40.271535,-121.01808700000001,1,19.85,0,0,None,4158,0,1,0,0,29,1,0.0,165.01000000000005,0.0,573.05,0,0,96137
1643,1,0,1,0,37,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,90.35,3419.3,0,56,22,6.99,3347,0,Carnelian Bay,1,1,Fiber Optic,39.227434,-120.091806,1,90.35,0,4,None,1943,1,0,1,1,37,1,75.22,258.63,0.0,3419.3,0,1,96140
1644,0,0,0,0,34,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Mailed check,109.8,3587.25,1,23,84,7.99,3410,1,San Diego,1,0,Fiber Optic,32.957195,-117.202542,0,114.192,0,0,None,28201,0,0,0,1,34,2,0.0,271.66,0.0,3587.25,1,1,92130
1645,0,1,0,0,42,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.65,3541.35,1,79,19,9.53,4871,1,San Diego,0,0,Fiber Optic,32.957195,-117.202542,0,88.03600000000002,0,0,None,28201,0,0,0,0,42,3,673.0,400.26,0.0,3541.35,0,0,92130
1646,0,0,1,1,59,1,1,DSL,1,1,0,0,One year,0,Mailed check,65.5,3801.3,0,57,25,14.49,5631,0,Kings Beach,0,0,Cable,39.246654,-120.029273,1,65.5,0,6,None,4806,1,0,1,0,59,0,0.0,854.91,0.0,3801.3,0,1,96143
1647,1,0,1,1,11,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),79.5,868.5,1,61,21,13.33,3469,1,San Diego,0,1,Cable,32.957195,-117.202542,1,82.68,0,1,Offer D,28201,0,0,1,0,11,3,182.0,146.63,0.0,868.5,0,0,92130
1648,1,1,1,1,60,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,80.95,4859.1,0,71,11,18.23,6214,0,Olympic Valley,0,1,Cable,39.191796999999994,-120.212401,1,80.95,1,10,None,942,0,0,1,0,60,1,0.0,1093.8,49.53,4859.1,0,1,96146
1649,0,0,0,0,27,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,56.15,1439.35,0,29,53,1.31,3056,0,Tahoe Vista,0,0,Fiber Optic,39.241240000000005,-120.05476499999999,0,56.15,0,0,None,678,1,0,0,0,27,3,763.0,35.37000000000001,0.0,1439.35,1,0,96148
1650,0,0,0,0,1,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Mailed check,85.8,85.8,1,30,65,34.47,2850,1,San Diego,0,0,DSL,32.957195,-117.202542,0,89.23200000000001,0,0,Offer E,28201,0,0,0,1,1,3,0.0,34.47,0.0,85.8,0,1,92130
1651,1,1,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.1,79.1,1,65,18,42.3,5001,1,San Diego,0,1,DSL,32.957195,-117.202542,0,82.264,0,0,None,28201,0,1,0,0,1,2,0.0,42.3,0.0,79.1,0,1,92130
1652,1,0,1,0,17,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,34.4,592.75,0,36,10,0.0,4207,0,Los Angeles,1,1,Fiber Optic,33.973616,-118.24902,1,34.4,0,1,None,54492,0,0,1,0,17,0,59.0,0.0,0.0,592.75,0,0,90001
1653,1,0,1,0,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.75,1185.95,0,31,0,18.68,4927,0,Los Angeles,0,1,NA,33.949255,-118.246978,1,20.75,0,9,None,44586,0,0,1,0,58,0,0.0,1083.44,0.0,1185.95,0,0,90002
1654,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,18.8,18.8,0,29,0,43.57,5160,0,Los Angeles,0,1,NA,33.964131,-118.272783,1,18.8,0,9,None,58198,0,0,1,0,1,3,0.0,43.57,0.0,18.8,1,0,90003
1655,0,0,1,1,3,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.3,134.5,1,19,56,44.46,4903,1,Los Angeles,0,0,Cable,34.076259,-118.31071499999999,1,46.072,0,1,Offer E,67852,0,0,1,1,3,3,75.0,133.38,0.0,134.5,1,0,90004
1656,0,0,0,0,53,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Electronic check,90.8,4921.2,0,50,19,2.51,5249,0,Los Angeles,1,0,Fiber Optic,34.059281,-118.30742,0,90.8,0,0,None,43019,0,0,0,0,53,0,0.0,133.03,0.0,4921.2,0,1,90005
1657,1,0,0,0,35,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,25.6,901.25,0,21,0,39.84,2980,0,Los Angeles,0,1,NA,34.048013,-118.293953,0,25.6,0,0,None,62784,0,0,0,0,35,0,0.0,1394.4,0.0,901.25,1,0,90006
1658,1,0,1,1,50,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Credit card (automatic),105.95,5341.8,1,37,14,20.88,5536,1,Los Angeles,1,1,DSL,34.027337,-118.28515,1,110.18799999999999,0,0,None,45025,0,1,0,1,50,3,748.0,1044.0,0.0,5341.8,0,0,90007
1659,1,0,1,1,68,1,1,DSL,0,1,0,1,Two year,0,Credit card (automatic),70.8,4859.95,0,35,10,11.12,5540,0,Los Angeles,0,1,Fiber Optic,34.008293,-118.34676599999999,1,70.8,0,1,None,30852,1,1,1,1,68,1,0.0,756.16,0.0,4859.95,0,1,90008
1660,1,0,1,0,47,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,25.4,1139.2,0,20,0,10.07,3159,0,Los Angeles,0,1,NA,34.062125,-118.31570900000001,1,25.4,0,1,None,1957,0,0,1,0,47,2,0.0,473.29,0.0,1139.2,1,0,90010
1661,0,1,1,0,65,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),108.8,7082.45,0,69,9,48.53,5225,0,Los Angeles,1,0,DSL,34.007090000000005,-118.25868100000001,1,108.8,0,4,None,101215,0,0,1,0,65,0,0.0,3154.4500000000007,21.52,7082.45,0,1,90011
1662,1,0,0,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.75,324.6,1,32,6,31.14,3965,1,Los Angeles,0,1,Fiber Optic,34.065875,-118.23872800000001,0,72.54,0,0,Offer E,30596,0,3,0,0,5,1,19.0,155.7,0.0,324.6,0,0,90012
1663,1,0,1,0,51,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.65,4812.75,1,44,10,21.08,4747,1,Los Angeles,0,1,DSL,34.044639000000004,-118.24041299999999,1,98.436,0,1,None,9732,0,1,1,1,51,4,481.0,1075.08,0.0,4812.75,0,0,90013
1664,0,0,0,0,46,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),96.05,4399.5,1,57,9,6.18,2712,1,Los Angeles,0,0,Fiber Optic,34.043144,-118.251977,0,99.89200000000001,0,0,None,3524,0,0,0,1,46,2,396.0,284.28,0.0,4399.5,0,0,90014
1665,0,0,0,0,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.85,663.55,0,51,8,42.41,4834,0,Los Angeles,0,0,Fiber Optic,34.039224,-118.26629299999999,0,76.85,0,0,Offer E,15140,0,0,0,0,9,3,5.31,381.69,0.0,663.55,0,1,90015
1666,0,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.25,174.65,0,41,0,15.86,2653,0,Los Angeles,0,0,NA,34.028331,-118.35433799999998,0,20.25,0,0,Offer E,46984,0,0,0,0,8,1,0.0,126.88,0.0,174.65,0,0,90016
1667,1,0,0,0,14,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),24.8,321.7,0,40,0,33.5,4527,0,Los Angeles,0,1,NA,34.052842,-118.264495,0,24.8,0,0,None,20692,0,0,0,0,14,0,0.0,469.0,0.0,321.7,0,0,90017
1668,0,0,0,0,45,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,115.65,5125.5,0,26,30,33.73,3974,0,Los Angeles,1,0,DSL,34.028735,-118.31723600000001,0,115.65,0,0,None,47143,1,0,0,1,45,2,0.0,1517.85,0.0,5125.5,1,1,90018
1669,0,0,0,0,8,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.6,548.9,0,21,42,1.28,2142,0,Los Angeles,0,0,Fiber Optic,34.049841,-118.33846000000001,0,74.6,0,0,Offer E,67520,0,0,0,0,8,0,0.0,10.24,0.0,548.9,1,1,90019
1670,1,1,0,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.15,50.15,1,68,13,39.78,3438,1,San Diego,1,1,Cable,32.898613,-117.202937,0,52.156000000000006,0,0,Offer E,4258,0,0,0,0,1,2,0.0,39.78,0.0,50.15,0,0,92121
1671,1,0,1,1,66,1,0,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),103.15,7031.3,0,40,19,39.45,4663,0,Los Angeles,1,1,Fiber Optic,34.029043,-118.23950400000001,1,103.15,2,7,None,3012,0,1,1,1,66,2,133.59,2603.7000000000007,0.0,7031.3,0,1,90021
1672,1,0,1,1,72,1,1,DSL,1,1,0,0,Two year,0,Credit card (automatic),72.1,5016.65,0,39,18,42.55,4658,0,Los Angeles,1,1,DSL,34.02381,-118.156582,1,72.1,0,5,None,68701,1,0,1,0,72,0,903.0,3063.6,0.0,5016.65,0,0,90022
1673,0,0,1,0,41,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),113.6,4594.95,1,41,11,5.01,4963,1,Los Angeles,1,0,Fiber Optic,34.017697,-118.200577,1,118.144,0,1,None,47487,1,0,1,1,41,3,505.0,205.41,0.0,4594.95,0,0,90023
1674,0,0,1,1,23,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.1,611.45,0,47,0,35.86,2267,0,Los Angeles,0,0,NA,34.066303000000005,-118.435479,1,25.1,2,4,None,44150,0,0,1,0,23,0,0.0,824.78,0.0,611.45,0,0,90024
1675,0,0,0,0,29,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,78.9,2384.15,1,37,8,44.33,3249,1,Los Angeles,0,0,DSL,34.046174,-118.44633300000001,0,82.05600000000003,0,0,None,41175,0,0,0,0,29,2,0.0,1285.57,0.0,2384.15,0,1,90025
1676,0,0,0,0,4,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,80.15,319.85,0,27,73,6.5,2841,0,Los Angeles,0,0,Fiber Optic,34.078990999999995,-118.26380400000001,0,80.15,0,0,Offer E,73686,0,0,0,0,4,1,0.0,26.0,0.0,319.85,1,1,90026
1677,1,0,1,1,6,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.4,153.3,0,58,0,31.73,2882,0,Los Angeles,0,1,NA,34.127194,-118.295647,1,25.4,3,8,Offer E,48727,0,0,1,0,6,0,0.0,190.38,0.0,153.3,0,0,90027
1678,0,1,1,0,67,1,1,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),105.4,7035.6,0,70,25,2.67,5703,0,Los Angeles,1,0,Fiber Optic,34.099869,-118.326843,1,105.4,0,3,None,30568,1,0,1,0,67,0,1759.0,178.89,0.0,7035.6,0,0,90028
1679,1,1,0,1,7,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.75,344.2,0,72,17,41.14,3779,0,Los Angeles,0,1,DSL,34.089953,-118.294824,0,45.75,1,0,None,41713,0,0,0,0,7,0,0.0,287.98,29.0,344.2,0,1,90029
1680,1,0,1,1,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,24.45,1431.65,0,64,0,32.93,5623,0,Los Angeles,0,1,NA,34.085807,-118.206617,1,24.45,0,7,None,38415,0,0,1,0,56,3,0.0,1844.08,0.0,1431.65,0,0,90031
1681,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.0,1849.2,0,56,0,39.98,6126,0,Los Angeles,0,0,NA,34.078821000000005,-118.177576,1,25.0,0,7,None,46960,0,0,1,0,72,0,0.0,2878.56,0.0,1849.2,0,0,90032
1682,1,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Electronic check,85.25,6083.1,0,64,30,16.58,6275,0,Los Angeles,1,1,DSL,34.050197999999995,-118.21094599999999,1,85.25,0,9,None,49431,0,1,1,1,72,1,1825.0,1193.7599999999998,0.0,6083.1,0,0,90033
1683,1,0,1,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.6,426.65,0,60,0,34.04,4617,0,Los Angeles,0,1,NA,34.030578000000006,-118.39961299999999,1,19.6,3,10,None,58218,0,0,1,0,23,1,0.0,782.92,0.0,426.65,0,0,90034
1684,0,0,0,1,35,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.15,1655.35,0,52,19,38.82,5879,0,Los Angeles,0,0,Fiber Optic,34.051809000000006,-118.383843,0,50.15,1,0,None,27799,0,0,0,0,35,0,31.45,1358.7,0.0,1655.35,0,1,90035
1685,1,1,1,0,27,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.55,1943.9,0,71,16,30.49,2534,0,Los Angeles,0,1,DSL,34.070291,-118.34919099999999,1,70.55,0,0,Offer C,32901,0,0,0,0,27,2,0.0,823.2299999999998,29.99,1943.9,0,1,90036
1686,0,0,1,1,26,1,1,DSL,0,1,0,0,Month-to-month,1,Electronic check,60.05,1616.15,1,35,14,22.33,2039,1,Los Angeles,0,0,Cable,34.002642,-118.287596,1,62.452,0,1,None,56709,1,2,1,0,26,4,0.0,580.5799999999998,0.0,1616.15,0,1,90037
1687,1,0,1,1,12,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,26.4,314.95,0,54,0,45.15,3277,0,Los Angeles,0,1,NA,34.088017,-118.327168,1,26.4,0,5,None,32562,0,0,1,0,12,0,0.0,541.8,0.0,314.95,0,0,90038
1688,0,0,0,0,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.15,804.85,0,33,0,8.36,3915,0,Los Angeles,0,0,NA,34.110845,-118.25959499999999,0,20.15,0,0,None,29310,0,0,0,0,40,2,0.0,334.4,0.0,804.85,0,0,90039
1689,1,0,1,1,7,0,No phone service,DSL,1,1,1,1,Month-to-month,0,Mailed check,58.85,465.7,0,21,47,0.0,3332,0,Los Angeles,1,1,DSL,33.994524,-118.149953,1,58.85,2,9,Offer E,9805,0,0,1,1,7,1,219.0,0.0,0.0,465.7,1,0,90040
1690,1,0,1,1,70,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Credit card (automatic),97.55,6669.05,0,62,53,32.38,4551,0,Los Angeles,0,1,DSL,34.137412,-118.20760700000001,1,97.55,3,8,None,27866,0,0,1,0,70,2,353.46,2266.600000000001,0.0,6669.05,0,1,90041
1691,1,0,1,1,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.65,1161.75,0,31,0,21.98,6315,0,Los Angeles,0,1,NA,34.11572,-118.19275400000001,1,19.65,1,7,None,64672,0,0,1,0,60,1,0.0,1318.8,0.0,1161.75,0,0,90042
1692,1,0,1,1,39,0,No phone service,DSL,0,0,0,0,One year,1,Credit card (automatic),25.25,947.75,0,27,48,0.0,4259,0,Los Angeles,0,1,DSL,33.988543,-118.33408100000001,1,25.25,0,8,None,44764,0,0,1,0,39,0,0.0,0.0,0.0,947.75,1,1,90043
1693,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),114.45,8375.05,0,53,8,6.29,6274,0,Los Angeles,1,1,Cable,33.952714,-118.292061,1,114.45,0,5,None,87383,1,0,1,1,72,0,670.0,452.88,0.0,8375.05,0,0,90044
1694,0,0,0,0,1,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,34.7,34.7,1,31,9,0.0,4476,1,Los Angeles,0,0,Fiber Optic,33.954017,-118.402447,0,36.088,0,0,Offer E,39334,0,0,0,0,1,4,0.0,0.0,0.0,34.7,0,0,90045
1695,1,0,1,1,54,1,1,DSL,0,1,1,0,One year,1,Electronic check,70.7,3770,0,49,28,48.45,5276,0,Los Angeles,0,1,DSL,34.108455,-118.362081,1,70.7,0,3,None,49839,1,0,1,0,54,0,1056.0,2616.3,0.0,3770.0,0,0,90046
1696,1,0,0,0,3,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.3,264.8,1,46,23,14.28,4934,1,Los Angeles,0,1,Cable,33.958149,-118.30844099999999,0,88.712,0,0,Offer E,47107,0,1,0,1,3,3,61.0,42.84,0.0,264.8,0,0,90047
1697,0,0,1,1,63,1,0,DSL,1,1,1,0,Two year,0,Credit card (automatic),75.55,4707.85,0,58,30,6.33,4626,0,Los Angeles,1,0,DSL,34.072945000000004,-118.37267,1,75.55,0,7,None,21739,1,0,1,0,63,2,1412.0,398.79,0.0,4707.85,0,0,90048
1698,1,0,1,1,71,1,1,Fiber optic,0,1,0,0,Two year,1,Electronic check,84.8,6152.4,0,40,75,33.67,5952,0,Los Angeles,0,1,Fiber Optic,34.091829,-118.491244,1,84.8,3,9,None,33523,1,0,1,0,71,1,461.43,2390.57,0.0,6152.4,0,1,90049
1699,0,0,0,0,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.65,958.1,0,56,0,23.25,5956,0,Los Angeles,0,0,NA,33.987945,-118.370442,0,20.65,0,0,None,8115,0,0,0,0,42,0,0.0,976.5,0.0,958.1,0,0,90056
1700,1,0,0,0,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.45,943,0,27,0,6.61,4342,0,Los Angeles,0,1,NA,34.061918,-118.27793899999999,0,20.45,0,0,None,44004,0,0,0,0,47,3,0.0,310.67,0.0,943.0,1,0,90057
1701,0,0,1,1,66,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),102.45,6615.15,1,41,13,48.77,4688,1,Los Angeles,1,0,Cable,34.001616999999996,-118.222274,1,106.54799999999999,0,1,Offer A,3642,0,4,1,1,66,2,0.0,3218.82,0.0,6615.15,0,1,90058
1702,0,0,1,0,21,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),104.4,2200.25,1,22,65,38.52,5570,1,Los Angeles,1,0,Cable,33.927254,-118.249826,1,108.576,0,1,Offer D,38128,0,0,1,1,21,4,0.0,808.9200000000002,0.0,2200.25,1,1,90059
1703,1,0,0,0,11,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,35.65,425.1,0,20,73,0.0,4986,0,Los Angeles,0,1,Fiber Optic,33.921279999999996,-118.27418600000001,0,35.65,0,0,None,24511,1,1,0,0,11,1,31.03,0.0,0.0,425.1,1,1,90061
1704,1,0,0,1,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.75,99.75,1,59,28,40.71,4214,1,Los Angeles,1,1,Cable,34.003553000000004,-118.30893300000001,0,103.74,0,0,None,29299,0,1,0,1,1,3,0.0,40.71,0.0,99.75,0,0,90062
1705,0,1,1,0,55,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,90.45,5044.8,0,68,21,22.74,5140,0,Los Angeles,1,0,Fiber Optic,34.044271,-118.18523700000001,1,90.45,0,4,None,55668,1,0,1,0,55,0,1059.0,1250.6999999999996,12.48,5044.8,0,0,90063
1706,1,0,0,0,69,1,1,Fiber optic,0,1,1,0,Two year,1,Credit card (automatic),97.65,6743.55,0,41,30,49.35,5709,0,Los Angeles,1,1,DSL,34.037251,-118.423573,0,97.65,0,0,Offer A,24505,1,0,0,0,69,0,0.0,3405.15,0.0,6743.55,0,1,90064
1707,0,1,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,73.85,196.4,0,74,25,46.65,2868,0,Los Angeles,1,0,Fiber Optic,34.108833000000004,-118.22971499999998,0,73.85,0,0,None,47534,0,0,0,0,3,2,0.0,139.95,0.0,196.4,0,1,90065
1708,1,0,0,0,4,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,74.4,299.7,1,39,3,28.89,3633,1,Los Angeles,1,1,Cable,34.002028,-118.430656,0,77.376,0,0,None,55204,1,0,0,1,4,4,9.0,115.56,0.0,299.7,0,0,90066
1709,1,1,0,0,30,1,1,DSL,0,0,1,0,Two year,1,Credit card (automatic),69.1,2093.9,0,69,30,19.92,3415,0,Los Angeles,1,1,Cable,34.057496,-118.413959,0,69.1,0,0,None,2527,1,0,0,0,30,0,0.0,597.6,21.08,2093.9,0,1,90067
1710,0,0,0,0,5,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,82.75,417.75,0,21,42,29.74,5269,0,Los Angeles,1,0,DSL,34.137411,-118.328915,0,82.75,0,0,Offer E,21728,1,0,0,0,5,1,0.0,148.7,0.0,417.75,1,1,90068
1711,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.4,1725.4,0,19,0,24.72,4412,0,West Hollywood,0,0,NA,34.093781,-118.38106100000002,1,24.4,0,1,Offer A,20408,0,0,1,0,71,2,0.0,1755.12,0.0,1725.4,1,0,90069
1712,0,0,0,0,29,1,1,DSL,0,1,0,0,One year,1,Electronic check,55.25,1620.2,0,28,69,39.35,5481,0,Los Angeles,0,0,Fiber Optic,34.052917,-118.255178,0,55.25,0,0,None,21,0,0,0,0,29,4,1118.0,1141.15,0.0,1620.2,1,0,90071
1713,1,0,1,0,52,1,1,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),61.35,3169.55,0,39,3,44.65,4729,0,Los Angeles,0,1,Cable,34.102084000000005,-118.451629,1,61.35,0,3,None,10470,1,1,1,0,52,1,0.0,2321.8,0.0,3169.55,0,1,90077
1714,1,0,0,0,68,1,1,DSL,1,1,0,1,One year,0,Credit card (automatic),76.75,5233.25,0,40,29,20.29,5395,0,Bell,1,1,Fiber Optic,33.970343,-118.17136799999999,0,76.75,0,0,Offer A,105285,0,0,0,1,68,2,151.76,1379.72,0.0,5233.25,0,1,90201
1715,0,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.4,967.85,0,61,0,47.5,2320,0,Beverly Hills,0,0,NA,34.099891,-118.41433799999999,1,19.4,1,9,None,21397,0,0,1,0,46,0,0.0,2185.0,0.0,967.85,0,0,90210
1716,1,0,0,0,8,1,0,DSL,0,0,0,1,Month-to-month,1,Credit card (automatic),54.75,438.05,0,63,26,30.53,5317,0,Beverly Hills,0,1,DSL,34.063947,-118.38300100000001,0,54.75,0,0,None,8321,0,0,0,1,8,1,11.39,244.24,0.0,438.05,0,1,90211
1717,1,0,1,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.7,1421.9,0,23,0,27.97,6436,0,Beverly Hills,0,1,NA,34.062095,-118.401508,1,19.7,0,10,Offer A,11355,0,0,1,0,72,0,0.0,2013.84,0.0,1421.9,1,0,90212
1718,0,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.9,323.15,0,38,0,25.62,2093,0,Compton,0,0,NA,33.88151,-118.234451,0,19.9,0,0,None,47305,0,0,0,0,17,0,0.0,435.54,0.0,323.15,0,0,90220
1719,1,0,0,0,3,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,107.95,318.6,0,42,28,12.66,5653,0,Compton,1,1,Cable,33.885811,-118.20645900000001,0,107.95,0,0,Offer E,51387,1,0,0,1,3,1,0.0,37.98,0.0,318.6,0,1,90221
1720,0,1,0,0,2,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),83.8,163.7,0,76,14,32.98,2885,0,Compton,0,0,Fiber Optic,33.912246,-118.236773,0,83.8,0,0,None,29825,0,0,0,0,2,1,0.0,65.96,0.0,163.7,0,1,90222
1721,0,0,0,0,9,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),74.25,639.65,1,23,84,13.86,5393,1,Culver City,0,0,DSL,33.993990999999994,-118.39703999999999,0,77.22,0,0,None,31963,0,1,0,1,9,5,537.0,124.74,0.0,639.65,1,0,90230
1722,0,0,0,0,51,0,No phone service,DSL,0,1,1,1,One year,1,Credit card (automatic),56.4,2928.5,0,52,24,0.0,4380,0,Culver City,1,0,DSL,34.019323,-118.391902,0,56.4,0,0,None,15195,0,0,0,1,51,0,703.0,0.0,0.0,2928.5,0,0,90232
1723,0,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.1,100.35,0,52,0,25.05,5874,0,Downey,0,0,NA,33.956228,-118.120993,1,20.1,1,4,Offer E,24908,0,0,1,0,6,1,0.0,150.3,0.0,100.35,0,0,90240
1724,0,0,1,0,3,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,94.9,273.2,0,51,7,2.97,2330,0,Downey,0,0,DSL,33.940884000000004,-118.128628,1,94.9,0,5,None,40152,0,0,1,1,3,1,19.0,8.91,0.0,273.2,0,0,90241
1725,0,1,0,0,17,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.2,1608.15,0,79,11,32.19,4425,0,Downey,0,0,Cable,33.921793,-118.140588,0,94.2,0,0,None,42459,0,0,0,1,17,1,0.0,547.23,36.4,1608.15,0,1,90242
1726,1,0,1,0,30,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,49.9,1441.95,0,62,8,5.56,3712,0,El Segundo,0,1,DSL,33.917145,-118.401554,1,49.9,0,4,None,16041,0,0,1,0,30,2,115.0,166.79999999999995,0.0,1441.95,0,0,90245
1727,1,0,0,0,31,1,1,DSL,0,1,1,0,Month-to-month,1,Electronic check,71.05,2168.15,0,39,24,6.4,4443,0,Gardena,0,1,DSL,33.890853,-118.29796699999999,0,71.05,0,0,None,47758,1,0,0,0,31,1,0.0,198.4,0.0,2168.15,0,1,90247
1728,0,0,0,0,45,1,0,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),81.65,3618.7,0,57,30,37.39,5937,0,Gardena,1,0,Cable,33.876482,-118.284077,0,81.65,0,0,Offer B,9960,1,0,0,1,45,1,0.0,1682.55,0.0,3618.7,0,1,90248
1729,1,0,1,0,64,1,1,Fiber optic,1,1,0,0,One year,0,Bank transfer (automatic),89.45,5692.65,0,30,48,13.8,5519,0,Gardena,1,1,Fiber Optic,33.90139,-118.315697,1,89.45,0,5,Offer B,26442,0,0,1,0,64,0,0.0,883.2,0.0,5692.65,0,1,90249
1730,1,0,0,0,1,1,1,DSL,0,0,1,0,Month-to-month,1,Electronic check,59.85,59.85,1,50,31,22.05,4017,1,Hawthorne,0,1,Cable,33.914775,-118.348083,0,62.24400000000001,0,0,None,93315,0,1,0,0,1,6,0.0,22.05,0.0,59.85,0,0,90250
1731,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.6,69.6,1,72,16,34.51,3438,1,Hermosa Beach,0,0,Cable,33.865320000000004,-118.396336,0,72.384,0,0,Offer E,18693,0,4,0,0,1,1,0.0,34.51,0.0,69.6,0,1,90254
1732,1,1,1,1,61,1,1,Fiber optic,0,1,1,1,One year,0,Electronic check,99.0,5969.3,0,80,22,4.51,5177,0,Huntington Park,0,1,Fiber Optic,33.97803,-118.217141,1,99.0,2,10,None,78114,0,1,1,1,61,2,0.0,275.11,21.17,5969.3,0,1,90255
1733,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.05,19.05,0,46,0,5.02,5279,0,Lawndale,0,1,NA,33.88856,-118.35181299999999,0,19.05,0,0,None,33300,0,0,0,0,1,0,0.0,5.02,0.0,19.05,0,0,90260
1734,1,0,0,0,9,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,45.4,418.8,1,54,22,0.0,5028,1,Lynwood,0,1,Fiber Optic,33.923573,-118.20066899999999,0,47.216,0,0,None,69850,0,2,0,1,9,4,92.0,0.0,0.0,418.8,0,0,90262
1735,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),114.45,8100.55,0,51,13,24.95,4700,0,Malibu,1,1,Fiber Optic,34.037037,-118.705803,1,114.45,1,0,Offer A,11,1,0,0,1,72,0,0.0,1796.4,0.0,8100.55,0,1,90263
1736,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.5,19.5,1,54,0,32.45,5211,1,Malibu,0,0,NA,34.074571999999996,-118.831181,0,19.5,0,0,None,19630,0,0,0,0,1,1,0.0,32.45,0.0,19.5,0,0,90265
1737,0,0,1,0,7,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.25,313.45,0,61,24,31.43,5014,0,Manhattan Beach,0,0,Cable,33.889632,-118.39737,1,44.25,0,4,None,33758,0,0,1,0,7,1,0.0,220.01,0.0,313.45,0,1,90266
1738,0,0,1,0,66,1,1,Fiber optic,0,1,0,0,One year,1,Bank transfer (automatic),90.55,6130.95,0,43,20,11.72,4958,0,Maywood,1,0,Fiber Optic,33.988572,-118.18656499999999,1,90.55,0,6,Offer A,28094,1,1,1,0,66,2,0.0,773.5200000000002,0.0,6130.95,0,1,90270
1739,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.9,69.9,1,56,13,45.5,3349,1,Pacific Palisades,0,1,DSL,34.079449,-118.54830600000001,0,72.69600000000001,0,0,None,22548,0,0,0,0,1,2,0.0,45.5,0.0,69.9,0,1,90272
1740,1,0,1,1,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.4,745.3,0,61,0,1.89,5918,0,Palos Verdes Peninsula,0,1,NA,33.788208000000004,-118.404955,1,20.4,1,2,Offer B,24979,0,0,1,0,40,2,0.0,75.6,0.0,745.3,0,0,90274
1741,1,0,0,0,16,1,1,DSL,0,1,0,1,Month-to-month,1,Bank transfer (automatic),71.4,1212.1,0,24,48,25.71,3360,0,Rancho Palos Verdes,1,1,Fiber Optic,33.753146,-118.36745900000001,0,71.4,0,0,None,41263,0,0,0,1,16,3,582.0,411.36,0.0,1212.1,1,0,90275
1742,0,0,0,0,2,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),87.15,183.75,1,50,7,6.2,4149,1,Redondo Beach,0,0,DSL,33.830453000000006,-118.384565,0,90.636,0,0,None,34191,0,0,0,0,2,3,13.0,12.4,0.0,183.75,0,0,90277
1743,1,0,1,0,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.85,1583.5,0,19,0,3.28,4833,0,Redondo Beach,0,1,NA,33.873395,-118.37019,1,24.85,0,9,Offer A,37322,0,0,1,0,67,2,0.0,219.76,0.0,1583.5,1,0,90278
1744,0,0,1,0,41,1,0,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),104.45,4162.05,0,45,14,9.85,2719,0,South Gate,1,0,Cable,33.944624,-118.19261499999999,1,104.45,0,2,Offer B,96267,0,0,1,1,41,1,0.0,403.85,0.0,4162.05,0,1,90280
1745,0,0,1,1,56,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.8,1119.9,0,58,0,48.56,4681,0,Topanga,0,0,NA,34.115192,-118.61017,1,19.8,1,2,Offer B,5451,0,0,1,0,56,0,0.0,2719.36,0.0,1119.9,0,0,90290
1746,0,0,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),116.45,8013.55,0,25,51,48.52,5567,0,Venice,1,0,DSL,33.991782,-118.479229,0,116.45,0,0,Offer A,31021,1,0,0,1,72,0,0.0,3493.44,0.0,8013.55,1,1,90291
1747,0,0,1,1,3,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),84.75,264.85,1,47,33,38.09,2014,1,Marina Del Rey,0,0,DSL,33.977468,-118.445475,1,88.14,0,1,None,18058,0,2,1,1,3,2,87.0,114.27,0.0,264.85,0,0,90292
1748,0,0,1,0,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.05,1102.4,0,58,0,32.72,4212,0,Playa Del Rey,0,0,NA,33.947305,-118.43984099999999,1,20.05,0,1,Offer B,11264,0,0,1,0,54,1,0.0,1766.88,0.0,1102.4,0,0,90293
1749,1,1,0,0,52,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,110.75,5832,0,75,25,23.04,4993,0,Inglewood,1,1,Fiber Optic,33.956445,-118.35863400000001,0,110.75,0,0,None,37527,1,0,0,1,52,0,0.0,1198.08,6.26,5832.0,0,1,90301
1750,0,0,0,0,50,1,0,Fiber optic,0,0,0,1,Two year,1,Bank transfer (automatic),89.7,4304.5,0,63,26,29.8,5306,0,Inglewood,1,0,Fiber Optic,33.975332,-118.35525200000001,0,89.7,0,0,Offer B,30779,1,1,0,1,50,2,1119.0,1490.0,0.0,4304.5,0,0,90302
1751,1,0,0,0,14,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,89.95,1178.4,1,40,30,28.65,5463,1,Inglewood,0,1,Cable,33.936291,-118.33263899999999,0,93.54799999999999,0,0,Offer D,27778,1,0,0,0,14,5,354.0,401.1,0.0,1178.4,0,0,90303
1752,1,0,1,0,27,1,0,DSL,1,0,0,0,One year,0,Credit card (automatic),48.7,1421.75,0,33,5,9.01,3560,0,Inglewood,0,1,Fiber Optic,33.936827,-118.359824,1,48.7,0,10,None,28680,0,0,1,0,27,2,0.0,243.27,0.0,1421.75,0,1,90304
1753,0,1,1,0,72,1,1,Fiber optic,1,1,0,0,Two year,1,Bank transfer (automatic),96.6,6827.5,0,70,20,28.09,5153,0,Inglewood,1,0,Fiber Optic,33.958134,-118.330905,1,96.6,0,10,None,13779,1,0,1,0,72,3,0.0,2022.48,0.0,6827.5,0,1,90305
1754,1,0,0,0,62,1,0,DSL,1,1,1,1,One year,1,Credit card (automatic),74.3,4698.05,0,56,30,38.33,5974,0,Santa Monica,0,1,Cable,34.015481,-118.49323100000001,0,74.3,0,0,Offer B,5221,0,0,0,1,62,0,1409.0,2376.46,0.0,4698.05,0,0,90401
1755,0,0,0,0,12,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,54.3,654.5,0,59,26,37.63,3854,0,Santa Monica,0,0,Fiber Optic,34.035849,-118.50350800000001,0,54.3,0,0,Offer D,11509,1,0,0,0,12,1,0.0,451.56000000000006,0.0,654.5,0,1,90402
1756,0,1,0,0,44,1,0,DSL,0,0,1,1,One year,0,Bank transfer (automatic),74.85,3268.05,0,76,17,7.72,3253,0,Santa Monica,1,0,DSL,34.031529,-118.491156,0,74.85,0,0,None,23559,1,0,0,1,44,2,0.0,339.68,17.91,3268.05,0,1,90403
1757,1,0,1,1,54,1,0,Fiber optic,0,1,0,0,Two year,1,Bank transfer (automatic),79.95,4362.05,0,31,75,46.7,4387,0,Santa Monica,0,1,DSL,34.026334000000006,-118.474222,1,79.95,8,2,Offer B,19975,1,0,1,0,54,3,0.0,2521.8,0.0,4362.05,0,1,90404
1758,0,0,0,0,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.05,1386.9,0,49,0,2.83,5740,0,Santa Monica,0,0,NA,34.005439,-118.477507,0,20.05,0,0,Offer A,26099,0,0,0,0,68,1,0.0,192.44,0.0,1386.9,0,0,90405
1759,1,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.4,415.4,0,20,0,31.02,4958,0,Torrance,0,1,NA,33.833698999999996,-118.31438700000001,0,19.4,0,0,Offer D,40705,0,0,0,0,20,1,0.0,620.4,0.0,415.4,1,0,90501
1760,1,0,1,1,50,1,1,DSL,0,0,0,0,One year,0,Bank transfer (automatic),54.9,2614.1,0,46,6,10.33,4322,0,Torrance,1,1,Fiber Optic,33.833181,-118.29206200000002,1,54.9,0,4,Offer B,17058,0,0,1,0,50,0,157.0,516.5,0.0,2614.1,0,0,90502
1761,1,0,0,0,58,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.45,1513.6,0,42,0,2.38,6490,0,Torrance,0,1,NA,33.840399,-118.353714,0,24.45,0,0,Offer B,41979,0,0,0,0,58,2,0.0,138.04,0.0,1513.6,0,0,90503
1762,1,0,1,1,35,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),89.65,3161.6,0,41,53,48.08,2622,0,Torrance,0,1,Fiber Optic,33.867257,-118.330794,1,89.65,3,4,None,31678,0,0,1,0,35,3,1676.0,1682.8,0.0,3161.6,0,0,90504
1763,0,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.4,80.95,0,31,13,10.81,4964,0,Torrance,0,0,Cable,33.807882,-118.34795700000001,0,45.4,0,0,None,34873,0,0,0,0,2,0,0.0,21.62,0.0,80.95,0,1,90505
1764,1,0,1,1,63,1,1,DSL,1,0,0,1,Two year,0,Mailed check,75.7,4676.7,0,35,21,12.15,5113,0,Whittier,1,1,DSL,34.007353,-118.03368300000001,1,75.7,0,3,Offer B,32050,1,0,1,1,63,1,982.0,765.45,0.0,4676.7,0,0,90601
1765,0,0,1,0,58,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),110.65,6526.65,0,35,18,37.95,4761,0,Whittier,1,0,Fiber Optic,33.972119,-118.02018799999999,1,110.65,0,8,Offer B,26265,0,0,1,1,58,1,0.0,2201.100000000001,0.0,6526.65,0,1,90602
1766,0,0,1,1,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.55,583.3,0,37,0,20.96,2269,0,Whittier,0,0,NA,33.945318,-117.992066,1,20.55,0,10,None,19109,0,0,1,0,27,0,0.0,565.9200000000002,0.0,583.3,0,0,90603
1767,0,0,1,0,71,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),115.15,8078.1,0,57,9,9.44,4144,0,Whittier,1,0,Cable,33.929704,-118.01208000000001,1,115.15,0,7,Offer A,37887,1,1,1,1,71,2,727.0,670.24,0.0,8078.1,0,0,90604
1768,0,0,0,0,63,1,0,DSL,0,0,0,1,One year,0,Credit card (automatic),58.55,3503.5,0,35,9,27.38,6312,0,Whittier,1,0,DSL,33.960891,-118.03222199999999,0,58.55,0,0,Offer B,38181,0,1,0,1,63,1,31.53,1724.9399999999996,0.0,3503.5,0,1,90605
1769,1,0,1,0,71,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),93.25,6669.45,0,40,7,26.56,6035,0,Whittier,1,1,DSL,33.976678,-118.065875,1,93.25,0,8,Offer A,32148,0,0,1,1,71,1,467.0,1885.76,0.0,6669.45,0,0,90606
1770,0,1,0,0,41,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,113.2,4689.5,1,66,25,27.95,3380,1,Buena Park,1,0,Cable,33.845706,-118.012204,0,117.728,0,0,None,44442,0,0,0,1,41,2,1172.0,1145.95,0.0,4689.5,0,0,90620
1771,1,1,0,0,13,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.5,1201.15,1,68,4,26.11,5394,1,Buena Park,0,1,Cable,33.874224,-117.99336799999999,0,94.12,0,0,None,33528,0,3,0,1,13,1,48.0,339.43,29.84,1201.15,0,0,90621
1772,1,0,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,79.0,143.65,1,33,23,48.66,5239,1,La Palma,0,1,Cable,33.850504,-118.039892,0,82.16,0,0,None,15505,0,2,0,0,2,2,33.0,97.32,0.0,143.65,0,0,90623
1773,0,0,1,1,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.35,1292.65,0,51,0,46.61,6303,0,Cypress,0,0,NA,33.818477,-118.038307,1,19.35,1,10,Offer A,47344,0,0,1,0,68,0,0.0,3169.48,0.0,1292.65,0,0,90630
1774,1,0,1,1,1,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,48.75,48.75,0,32,22,26.26,5068,0,La Habra,0,1,Cable,33.940619,-117.9513,1,48.75,2,10,None,67354,0,1,1,0,1,4,0.0,26.26,0.0,48.75,0,0,90631
1775,1,1,0,0,65,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,109.05,7108.2,0,67,10,4.4,5692,0,La Mirada,1,1,DSL,33.902045,-118.00896100000001,0,109.05,0,0,None,47568,1,0,0,1,65,1,0.0,286.0,34.67,7108.2,0,1,90638
1776,1,1,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.0,1802.55,0,77,0,28.99,4055,0,Montebello,0,1,NA,34.015217,-118.10996200000001,1,25.0,0,0,None,62425,0,0,0,0,72,1,0.0,2087.28,28.93,1802.55,0,0,90640
1777,0,0,0,0,28,1,1,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),54.9,1505.15,0,37,11,3.25,2885,0,Norwalk,0,0,Fiber Optic,33.905963,-118.08263000000001,0,54.9,0,0,None,103214,1,0,0,0,28,1,0.0,91.0,0.0,1505.15,0,1,90650
1778,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.75,1859.1,0,54,0,47.69,4185,0,Pico Rivera,0,1,NA,33.989523999999996,-118.089299,1,24.75,2,3,Offer A,63288,0,0,1,0,72,1,0.0,3433.68,0.0,1859.1,0,0,90660
1779,0,0,0,0,2,1,0,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,91.15,168.5,0,36,12,46.78,2686,0,Santa Fe Springs,0,0,DSL,33.933565,-118.062611,0,91.15,0,0,None,16271,0,0,0,0,2,0,20.0,93.56,0.0,168.5,0,0,90670
1780,0,0,0,1,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.15,390.85,1,39,0,8.95,4931,1,Stanton,0,0,NA,33.801869,-117.99506799999999,0,20.15,0,0,Offer D,29694,0,0,0,0,18,1,0.0,161.1,0.0,390.85,0,0,90680
1781,1,1,1,0,60,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,104.35,6339.45,0,80,15,22.95,4040,0,Artesia,1,1,Fiber Optic,33.867593,-118.08063700000001,1,104.35,0,2,None,16398,0,0,1,1,60,1,951.0,1377.0,41.23,6339.45,0,0,90701
1782,0,1,0,0,26,1,1,DSL,0,0,0,1,Month-to-month,1,Electronic check,66.05,1652.4,0,79,15,12.09,3225,0,Cerritos,0,0,Cable,33.8681,-118.067402,0,66.05,0,0,None,51556,1,0,0,1,26,1,248.0,314.34,47.73,1652.4,0,0,90703
1783,1,0,0,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.65,71.65,1,60,18,17.54,2377,1,Avalon,0,1,DSL,33.391181,-118.421305,0,74.516,0,0,None,3699,0,2,0,0,1,3,0.0,17.54,0.0,71.65,0,0,90704
1784,0,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,77.5,1,35,0,37.66,5984,1,Bellflower,0,0,NA,33.887676,-118.12728899999999,0,20.35,0,0,None,72893,0,0,0,0,4,1,0.0,150.64,0.0,77.5,0,0,90706
1785,1,0,1,1,68,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),92.2,6392.85,0,39,20,38.38,4451,0,Harbor City,1,1,Cable,33.798266,-118.30023700000001,1,92.2,0,4,Offer A,24660,1,0,1,1,68,2,1279.0,2609.84,0.0,6392.85,0,0,90710
1786,0,0,0,0,38,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),84.25,3264.5,1,26,45,17.66,2885,1,Lakewood,1,0,DSL,33.840524,-118.148403,0,87.62,0,0,None,30173,1,0,0,1,38,2,1469.0,671.08,0.0,3264.5,1,0,90712
1787,0,1,1,0,42,1,1,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),105.2,4599.15,0,79,7,35.38,5573,0,Lakewood,1,0,Cable,33.847755,-118.112532,1,105.2,0,2,None,27563,0,0,1,1,42,1,322.0,1485.96,40.46,4599.15,0,0,90713
1788,0,0,1,0,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.6,1134.25,0,54,0,23.28,6064,0,Lakewood,0,0,NA,33.841027000000004,-118.078097,1,19.6,0,10,Offer B,20890,0,0,1,0,57,0,0.0,1326.96,0.0,1134.25,0,0,90715
1789,1,0,1,0,54,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,30.4,1621.35,0,45,9,0.0,4778,0,Hawaiian Gardens,0,1,Fiber Optic,33.830431,-118.07407099999999,1,30.4,0,9,Offer B,14852,0,0,1,0,54,1,146.0,0.0,0.0,1621.35,0,0,90716
1790,0,0,0,0,12,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Bank transfer (automatic),78.1,947.3,1,32,20,42.55,4741,1,Lomita,0,0,Fiber Optic,33.794209,-118.31735400000001,0,81.22399999999999,0,0,Offer D,21065,0,0,0,1,12,5,189.0,510.6,0.0,947.3,0,0,90717
1791,0,0,1,0,44,1,0,DSL,1,1,0,0,One year,1,Mailed check,61.5,2722.2,0,60,20,44.87,2059,0,Los Alamitos,1,0,Fiber Optic,33.794990000000006,-118.065591,1,61.5,0,8,Offer B,21343,0,0,1,0,44,2,0.0,1974.28,0.0,2722.2,0,1,90720
1792,1,0,1,1,42,1,1,DSL,1,1,1,0,Month-to-month,1,Bank transfer (automatic),69.4,3058.3,0,64,17,16.67,4701,0,Paramount,0,1,Fiber Optic,33.897121999999996,-118.164432,1,69.4,1,10,Offer B,55306,0,1,1,0,42,1,0.0,700.1400000000001,0.0,3058.3,0,1,90723
1793,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.75,1769.6,0,27,0,35.33,6232,0,San Pedro,0,1,NA,33.736387,-118.28436299999998,1,24.75,1,1,Offer A,58639,0,0,1,0,72,1,0.0,2543.76,0.0,1769.6,1,0,90731
1794,0,0,1,1,71,1,1,DSL,1,1,1,1,Two year,0,Mailed check,91.05,6293.75,0,26,76,9.5,4644,0,San Pedro,1,0,Fiber Optic,33.744119,-118.31448,1,91.05,0,3,Offer A,21279,1,0,1,1,71,0,0.0,674.5,0.0,6293.75,1,1,90732
1795,0,0,1,0,19,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Mailed check,89.65,1761.05,1,20,52,21.71,3046,1,Seal Beach,1,0,Cable,33.75462,-118.071128,1,93.236,0,1,Offer D,24180,0,1,1,1,19,2,916.0,412.49,0.0,1761.05,1,0,90740
1796,0,0,1,0,23,1,1,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),73.65,1642.75,0,20,48,14.53,2590,0,Sunset Beach,0,0,Cable,33.719221000000005,-118.073596,1,73.65,0,5,Offer D,1107,1,0,1,1,23,0,0.0,334.19,0.0,1642.75,1,1,90742
1797,0,0,0,0,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.4,578.5,0,35,0,9.27,3986,0,Surfside,0,0,NA,33.728273,-118.08530400000001,0,19.4,0,0,None,174,0,1,0,0,30,2,0.0,278.1,0.0,578.5,0,0,90743
1798,1,0,0,0,35,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),26.2,954.9,0,40,0,49.13,4419,0,Wilmington,0,1,NA,33.782068,-118.26226299999999,0,26.2,0,0,None,53323,0,0,0,0,35,2,0.0,1719.5500000000004,0.0,954.9,0,0,90744
1799,0,0,0,0,10,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,98.7,973.25,1,35,31,37.36,5561,1,Carson,0,0,Cable,33.822295000000004,-118.26411,0,102.648,0,0,Offer D,55486,0,0,0,1,10,4,302.0,373.6,0.0,973.25,0,0,90745
1800,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),43.85,43.85,0,54,27,15.9,5913,0,Carson,0,1,Fiber Optic,33.859171,-118.25227199999999,0,43.85,0,0,None,25566,0,0,0,0,1,1,0.0,15.9,0.0,43.85,0,0,90746
1801,1,0,0,0,22,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.7,1490.4,0,22,42,15.77,4838,0,Long Beach,0,1,Fiber Optic,33.752524,-118.21073700000001,0,69.7,0,0,Offer D,38427,0,1,0,0,22,2,626.0,346.94,0.0,1490.4,1,0,90802
1802,1,0,1,1,7,0,No phone service,DSL,1,1,0,0,Two year,0,Mailed check,38.55,280,0,26,58,0.0,3345,0,Long Beach,1,1,DSL,33.760458,-118.129725,1,38.55,0,5,None,31352,0,1,1,0,7,2,162.0,0.0,0.0,280.0,1,0,90803
1803,0,0,0,0,36,0,No phone service,DSL,1,1,0,1,Two year,1,Mailed check,53.1,1901.25,0,46,9,0.0,2751,0,Long Beach,1,0,Fiber Optic,33.783046999999996,-118.1486,0,53.1,0,0,None,43467,1,0,0,1,36,0,0.0,0.0,0.0,1901.25,0,1,90804
1804,0,0,1,1,34,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.65,716.4,0,39,0,9.66,5099,0,Long Beach,0,0,NA,33.864622,-118.179626,1,20.65,1,7,None,91664,0,1,1,0,34,1,0.0,328.44,0.0,716.4,0,0,90805
1805,1,0,1,1,72,1,1,DSL,1,1,0,0,Two year,0,Credit card (automatic),64.45,4720,0,25,48,32.67,6330,0,Long Beach,1,1,Fiber Optic,33.802664,-118.179971,1,64.45,0,1,Offer A,49647,0,0,1,0,72,0,2266.0,2352.24,0.0,4720.0,1,0,90806
1806,1,0,1,1,36,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.1,930.95,0,48,0,34.79,3040,0,Long Beach,0,1,NA,33.830099,-118.182239,1,25.1,1,9,None,31556,0,0,1,0,36,1,0.0,1252.44,0.0,930.95,0,0,90807
1807,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,76.35,76.35,1,63,10,7.26,5613,1,Long Beach,1,0,DSL,33.823943,-118.11133500000001,0,79.404,0,0,None,37417,0,0,0,0,1,5,0.0,7.26,0.0,76.35,0,0,90808
1808,0,0,0,0,23,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.15,1676.95,1,51,12,33.44,5216,1,Long Beach,0,0,Cable,33.819814,-118.222416,0,82.316,0,0,Offer D,35656,0,2,0,0,23,2,0.0,769.1199999999999,0.0,1676.95,0,1,90810
1809,1,1,1,0,32,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.0,2642.05,1,69,25,5.99,4584,1,Long Beach,0,1,DSL,33.781086,-118.199049,1,88.4,0,1,None,63136,0,2,1,1,32,3,661.0,191.68,49.57,2642.05,0,0,90813
1810,0,0,1,1,71,1,1,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),95.15,6770.85,0,35,19,34.53,5647,0,Long Beach,1,0,Fiber Optic,33.771612,-118.14386599999999,1,95.15,1,3,Offer A,19034,1,0,1,0,71,0,1286.0,2451.63,0.0,6770.85,0,0,90814
1811,0,1,0,0,23,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,79.35,1835.3,0,66,18,8.72,3558,0,Long Beach,1,0,Cable,33.797638,-118.11662,0,79.35,0,0,None,38902,0,0,0,0,23,0,33.04,200.56,15.41,1835.3,0,1,90815
1812,1,0,1,0,17,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),96.65,1588.25,0,33,5,28.83,5228,0,Long Beach,1,1,Fiber Optic,33.778436,-118.118648,1,96.65,0,1,Offer D,425,0,0,1,1,17,0,0.0,490.11,0.0,1588.25,0,1,90822
1813,1,0,0,0,1,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,75.5,75.5,0,26,52,5.63,2954,0,Altadena,1,1,DSL,34.196837,-118.14223600000001,0,75.5,0,0,None,36243,1,2,0,1,1,1,0.0,5.63,0.0,75.5,1,1,91001
1814,1,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.7,258.35,0,44,0,4.71,5104,0,Arcadia,0,1,NA,34.137319,-118.02983700000001,1,19.7,3,7,Offer D,30028,0,0,1,0,12,2,0.0,56.52,0.0,258.35,0,0,91006
1815,0,0,1,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.5,1502.25,0,51,0,43.91,6302,0,Arcadia,0,0,NA,34.128284,-118.04773200000001,1,20.5,0,6,Offer A,30933,0,1,1,0,72,1,0.0,3161.5199999999995,0.0,1502.25,0,0,91007
1816,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.2,19.2,0,33,0,35.88,4629,0,Duarte,0,1,NA,34.145695,-117.95982,0,19.2,0,0,None,27414,0,0,0,0,1,0,0.0,35.88,0.0,19.2,0,0,91010
1817,1,1,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,0,Bank transfer (automatic),98.35,6929.4,0,65,30,44.61,6120,0,La Canada Flintridge,0,1,DSL,34.234912,-118.153729,1,98.35,0,0,None,20200,0,0,0,1,72,0,0.0,3211.92,0.0,6929.4,0,1,91011
1818,1,0,1,1,60,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),74.35,4453.3,0,50,57,38.44,5100,0,Monrovia,0,1,Fiber Optic,34.1528,-118.000482,1,74.35,4,9,Offer B,41067,0,0,1,0,60,2,0.0,2306.4,0.0,4453.3,0,1,91016
1819,0,0,1,1,61,0,No phone service,DSL,0,1,1,0,Two year,0,Credit card (automatic),51.35,3244.4,0,38,17,0.0,4159,0,Montrose,1,0,Fiber Optic,34.2112,-118.230625,1,51.35,0,10,Offer B,7527,1,0,1,0,61,1,552.0,0.0,0.0,3244.4,0,0,91020
1820,0,0,1,0,6,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.65,323.45,0,27,27,5.69,4227,0,Sierra Madre,0,0,DSL,34.168686,-118.057505,1,45.65,0,9,Offer E,10558,0,0,1,0,6,0,87.0,34.14,0.0,323.45,1,0,91024
1821,1,1,1,0,32,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,85.3,2661.1,1,76,11,49.6,2712,1,South Pasadena,0,1,Cable,34.110444,-118.156957,1,88.712,0,1,None,23984,0,2,1,1,32,5,293.0,1587.2,0.0,2661.1,0,0,91030
1822,0,0,0,1,31,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),86.55,2697.4,1,44,30,33.38,4198,1,Sunland,0,0,Cable,34.282703999999995,-118.312929,0,90.012,0,0,None,18752,0,0,0,0,31,2,809.0,1034.78,0.0,2697.4,0,0,91040
1823,1,0,0,0,19,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),73.85,1424.5,1,47,15,1.79,2251,1,Tujunga,0,1,Cable,34.296574,-118.24483899999998,0,76.804,0,0,Offer D,26753,0,1,0,0,19,2,0.0,34.01,0.0,1424.5,0,1,91042
1824,1,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.3,1401.15,0,29,0,27.16,5265,0,Pasadena,0,1,NA,34.146634999999996,-118.139225,1,20.3,1,9,Offer A,16812,0,0,1,0,72,3,0.0,1955.52,0.0,1401.15,1,0,91101
1825,0,0,0,0,32,1,1,DSL,0,1,0,0,Month-to-month,1,Electronic check,54.2,1739.6,0,42,3,32.02,4454,0,Pasadena,0,0,DSL,34.167465,-118.165327,0,54.2,0,0,None,27891,0,0,0,0,32,0,0.0,1024.64,0.0,1739.6,0,1,91103
1826,1,0,1,0,65,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,90.65,5931,0,52,2,19.84,6358,0,Pasadena,0,1,Fiber Optic,34.165383,-118.123752,1,90.65,0,1,Offer B,38460,0,0,1,1,65,2,0.0,1289.6,0.0,5931.0,0,1,91104
1827,0,0,1,1,45,0,No phone service,DSL,1,0,1,1,Month-to-month,1,Bank transfer (automatic),50.9,2333.85,0,54,18,0.0,3937,0,Pasadena,0,0,Cable,34.13946,-118.16664899999999,1,50.9,2,10,Offer B,10253,0,0,1,1,45,0,420.0,0.0,0.0,2333.85,0,0,91105
1828,1,0,0,0,42,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,25.05,949.85,0,20,0,27.64,3756,0,Pasadena,0,1,NA,34.139402000000004,-118.128658,0,25.05,0,0,None,23742,0,0,0,0,42,0,0.0,1160.88,0.0,949.85,1,0,91106
1829,1,0,0,0,8,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.85,572.45,0,64,7,11.58,5514,0,Pasadena,0,1,DSL,34.159007,-118.08735300000001,0,74.85,0,0,Offer E,32369,0,0,0,0,8,0,40.0,92.64,0.0,572.45,0,0,91107
1830,1,0,0,1,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.5,696.8,0,38,0,16.94,3114,0,San Marino,0,1,NA,34.122671000000004,-118.11291100000001,0,20.5,2,0,None,13158,0,0,0,0,32,0,0.0,542.08,0.0,696.8,0,0,91108
1831,0,1,1,0,22,1,1,DSL,1,1,0,0,Month-to-month,1,Mailed check,63.55,1381.8,0,73,25,17.22,2136,0,Glendale,0,0,DSL,34.17051,-118.28946299999998,1,63.55,0,5,Offer D,23981,1,0,1,0,22,1,0.0,378.84,0.0,1381.8,0,1,91201
1832,1,1,1,0,57,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,44.85,2572.95,1,70,3,0.0,5172,1,Glendale,0,1,Cable,34.167926,-118.26753899999999,1,46.64400000000001,0,1,None,21990,0,0,1,1,57,7,77.0,0.0,12.07,2572.95,0,0,91202
1833,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,47.95,47.95,0,33,25,46.23,5092,0,Glendale,0,1,Fiber Optic,34.153338,-118.262974,0,47.95,0,0,Offer E,14493,0,1,0,0,1,2,0.0,46.23,0.0,47.95,0,0,91203
1834,1,1,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.1,45.1,1,71,15,15.28,4499,1,Glendale,0,1,Cable,34.136306,-118.26036,0,46.903999999999996,0,0,Offer E,17015,0,1,0,0,1,9,0.0,15.28,0.0,45.1,0,0,91204
1835,0,0,1,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.0,45,0,25,52,40.63,5669,0,Glendale,0,0,Cable,34.13658,-118.24583899999999,1,45.0,0,7,Offer E,41390,0,0,1,0,1,1,0.0,40.63,0.0,45.0,1,1,91205
1836,1,0,0,0,24,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.0,2122.45,1,44,2,24.76,3068,1,Glendale,0,1,Cable,34.162515,-118.203869,0,99.84,0,0,None,31297,1,2,0,1,24,2,42.0,594.24,0.0,2122.45,0,0,91206
1837,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.05,20.05,1,57,0,12.0,4710,1,Glendale,0,1,NA,34.182378,-118.262922,0,20.05,0,0,None,9864,0,1,0,0,1,3,0.0,12.0,0.0,20.05,0,0,91207
1838,1,1,0,0,54,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,90.05,4931.8,0,69,14,18.58,5232,0,Glendale,0,1,Fiber Optic,34.195386,-118.23850800000001,0,90.05,0,0,None,16910,0,0,0,0,54,1,0.0,1003.32,0.0,4931.8,0,1,91208
1839,0,0,0,0,4,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.3,116.95,0,24,0,9.75,3808,0,La Crescenta,0,0,NA,34.239636,-118.245259,0,25.3,0,0,Offer E,29110,0,0,0,0,4,1,0.0,39.0,0.0,116.95,1,0,91214
1840,1,0,1,1,65,1,1,Fiber optic,1,0,1,1,Two year,0,Bank transfer (automatic),108.65,6937.95,1,53,8,41.88,6120,1,Agoura Hills,1,1,DSL,34.129058,-118.75978799999999,1,112.996,0,0,None,25303,1,0,0,1,65,2,55.5,2722.2000000000007,0.0,6937.95,0,1,91301
1841,0,0,1,0,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,24.3,1261.7,0,23,0,21.21,5052,0,Calabasas,0,0,NA,34.130860999999996,-118.68346000000001,1,24.3,0,7,None,23661,0,0,1,0,56,2,0.0,1187.76,0.0,1261.7,1,0,91302
1842,1,0,0,0,45,1,0,DSL,1,0,1,1,Month-to-month,1,Electronic check,75.95,3273.8,0,61,6,10.36,2185,0,Canoga Park,1,1,Fiber Optic,34.19829,-118.602203,0,75.95,0,0,None,23519,0,1,0,1,45,1,0.0,466.2,0.0,3273.8,0,1,91303
1843,0,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.7,1415.85,0,22,0,22.36,5921,0,Canoga Park,0,0,NA,34.224377000000004,-118.63265600000001,1,19.7,2,5,None,49242,0,0,1,0,71,1,0.0,1587.56,0.0,1415.85,1,0,91304
1844,1,0,1,0,59,1,0,DSL,1,1,1,0,One year,0,Credit card (automatic),66.4,3958.2,0,49,4,16.06,6432,0,Winnetka,1,1,Fiber Optic,34.209532,-118.57756299999998,1,66.4,0,3,None,43857,0,0,1,0,59,1,158.0,947.54,0.0,3958.2,0,0,91306
1845,1,0,0,0,69,0,No phone service,DSL,0,1,0,0,One year,1,Bank transfer (automatic),35.75,2492.25,0,37,19,0.0,4043,0,West Hills,1,1,Fiber Optic,34.199787,-118.68493000000001,0,35.75,0,0,None,23637,0,0,0,0,69,1,0.0,0.0,0.0,2492.25,0,1,91307
1846,1,0,0,0,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,18.8,279.2,0,62,0,17.17,2916,0,Chatsworth,0,1,NA,34.294142,-118.60388300000001,0,18.8,0,0,Offer D,35325,0,0,0,0,19,2,0.0,326.23,0.0,279.2,0,0,91311
1847,0,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.4,1083,0,24,0,27.75,5366,0,Encino,0,0,NA,34.150354,-118.51829199999999,1,19.4,2,8,None,27614,0,0,1,0,55,1,0.0,1526.25,0.0,1083.0,1,0,91316
1848,0,0,0,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.3,755.5,0,48,0,32.63,4705,0,Newbury Park,0,0,NA,34.172071,-118.946262,0,19.3,0,0,None,37779,0,0,0,0,38,0,0.0,1239.94,0.0,755.5,0,0,91320
1849,1,0,0,0,10,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.55,402.6,1,28,76,34.44,4097,1,Newhall,0,1,Fiber Optic,34.370378,-118.50411799999999,0,47.372,0,0,Offer D,30742,0,0,0,1,10,3,0.0,344.4,0.0,402.6,1,1,91321
1850,0,1,1,0,47,1,1,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),67.45,3252,0,78,24,46.77,4074,0,Northridge,1,0,Fiber Optic,34.238208,-118.55028999999999,1,67.45,0,1,None,25751,0,0,1,0,47,2,78.05,2198.19,0.0,3252.0,0,1,91324
1851,0,0,1,0,2,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,35.1,68.75,1,36,13,0.0,2643,1,Northridge,0,0,Cable,34.236683,-118.51758799999999,1,36.50400000000001,0,1,Offer E,32307,0,0,1,1,2,1,0.0,0.0,0.0,68.75,0,1,91325
1852,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),46.2,46.2,1,47,23,48.58,4167,1,Porter Ranch,0,1,Fiber Optic,34.281911,-118.55621799999999,0,48.048,0,0,Offer E,28067,0,2,0,0,1,2,0.0,48.58,0.0,46.2,0,0,91326
1853,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.15,45.15,1,29,76,30.92,5828,1,Pacoima,0,0,Cable,34.255441999999995,-118.421314,0,46.956,0,0,Offer E,97318,0,0,0,1,1,3,0.0,30.92,0.0,45.15,1,0,91331
1854,1,1,0,0,1,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Electronic check,43.3,43.3,1,75,29,0.0,4972,1,Reseda,1,1,DSL,34.200175,-118.540958,0,45.032,0,0,Offer E,68018,0,0,0,0,1,1,0.0,0.0,0.0,43.3,0,1,91335
1855,1,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.1,936.85,0,35,0,14.91,3392,0,San Fernando,0,1,NA,34.286131,-118.435969,1,20.1,2,4,None,33389,0,1,1,0,46,1,0.0,685.86,0.0,936.85,0,0,91340
1856,0,1,0,0,38,1,0,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),57.15,2250.65,1,67,30,26.1,3110,1,Sylmar,0,0,Cable,34.321621,-118.399841,0,59.43600000000001,0,0,None,81986,0,1,0,0,38,3,67.52,991.8,0.0,2250.65,0,1,91342
1857,0,0,1,0,65,1,0,DSL,1,0,0,0,Two year,0,Credit card (automatic),58.9,3857.1,0,22,71,34.31,5657,0,North Hills,1,0,DSL,34.238802,-118.48229599999999,1,58.9,0,5,None,57017,1,0,1,0,65,2,0.0,2230.15,0.0,3857.1,1,1,91343
1858,0,0,1,0,19,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,73.2,1441.1,1,31,24,25.75,4718,1,Granada Hills,0,0,Cable,34.291273,-118.505104,1,76.128,0,1,Offer D,48867,0,0,1,0,19,5,346.0,489.25,0.0,1441.1,0,0,91344
1859,1,0,0,0,52,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,85.35,4338.6,1,46,13,48.13,6402,1,Mission Hills,0,1,Cable,34.266389000000004,-118.459744,0,88.764,0,0,None,17112,0,0,0,1,52,2,0.0,2502.76,0.0,4338.6,0,1,91345
1860,1,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.45,1378.45,0,21,0,11.3,5497,0,Santa Clarita,0,1,NA,34.502432,-118.41458999999999,1,19.45,3,6,None,40077,0,0,1,0,71,0,0.0,802.3000000000002,0.0,1378.45,1,0,91350
1861,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.95,45.95,1,23,33,5.12,4888,1,Canyon Country,0,0,Cable,34.422519,-118.420717,0,47.788,0,0,Offer E,59259,0,0,0,1,1,3,0.0,5.12,0.0,45.95,1,0,91351
1862,0,1,0,0,52,0,No phone service,DSL,0,1,1,0,Month-to-month,1,Electronic check,50.5,2566.3,0,78,23,0.0,5185,0,Sun Valley,1,0,Cable,34.231053,-118.338307,0,50.5,0,0,None,46639,1,0,0,0,52,0,0.0,0.0,0.0,2566.3,0,1,91352
1863,1,0,1,0,6,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,25.1,171,0,37,0,47.29,5161,0,Valencia,0,1,NA,34.457005,-118.57372600000001,1,25.1,0,4,None,17846,0,0,1,0,6,0,0.0,283.74,0.0,171.0,0,0,91354
1864,0,1,1,0,26,1,0,DSL,0,0,0,1,One year,0,Mailed check,60.7,1597.4,0,76,17,17.12,2502,0,Valencia,1,0,Fiber Optic,34.43987,-118.644609,1,60.7,0,2,None,24977,0,0,1,0,26,2,0.0,445.12,0.0,1597.4,0,1,91355
1865,1,1,0,0,48,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,99.0,4744.35,0,71,2,5.87,3061,0,Tarzana,0,1,DSL,34.157137,-118.548511,0,99.0,0,0,None,27424,0,0,0,0,48,1,0.0,281.76,0.0,4744.35,0,1,91356
1866,0,0,1,1,64,1,1,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),104.4,6721.6,0,42,11,13.95,5133,0,Thousand Oaks,0,0,Fiber Optic,34.214054,-118.88108999999999,1,104.4,2,4,None,42526,1,1,1,1,64,1,739.0,892.8,0.0,6721.6,0,0,91360
1867,0,0,0,0,3,1,0,Fiber optic,0,1,1,0,Month-to-month,0,Electronic check,83.75,247.25,1,55,4,46.36,4852,1,Westlake Village,0,0,DSL,34.130992,-118.894673,0,87.10000000000002,0,0,Offer E,18735,0,0,0,0,3,7,0.0,139.07999999999998,0.0,247.25,0,1,91361
1868,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),44.05,44.05,0,49,10,30.73,5925,0,Thousand Oaks,0,1,Cable,34.191842,-118.822796,0,44.05,0,0,Offer E,33057,0,0,0,0,1,2,0.0,30.73,0.0,44.05,0,1,91362
1869,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.1,1734.65,0,48,0,19.64,4264,0,Woodland Hills,0,1,NA,34.153733,-118.59340800000001,1,24.1,1,0,None,25988,0,0,0,0,72,2,0.0,1414.08,0.0,1734.65,0,0,91364
1870,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.55,45.55,0,50,4,16.34,3173,0,Woodland Hills,0,1,Fiber Optic,34.178067999999996,-118.61571399999998,0,45.55,0,0,Offer E,36123,0,0,0,0,1,0,0.0,16.34,0.0,45.55,0,0,91367
1871,0,0,1,1,51,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,93.8,4539.35,0,41,75,27.23,5457,0,Oak Park,0,0,Fiber Optic,34.19225,-118.77687399999999,1,93.8,3,9,None,14814,0,0,1,1,51,1,340.45,1388.73,0.0,4539.35,0,1,91377
1872,0,0,1,1,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.7,804.25,0,45,0,23.95,2902,0,Stevenson Ranch,0,0,NA,34.364153,-118.615583,1,19.7,1,1,None,9937,0,2,1,0,41,1,0.0,981.95,0.0,804.25,0,0,91381
1873,0,0,1,1,72,1,0,DSL,1,1,1,0,Two year,1,Credit card (automatic),70.65,5011.15,0,59,22,43.12,5176,0,Castaic,1,0,Cable,34.506627,-118.699048,1,70.65,0,6,None,22177,0,0,1,0,72,2,1102.0,3104.64,0.0,5011.15,0,0,91384
1874,0,0,1,0,43,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),86.45,3574.5,0,64,14,21.08,3110,0,Van Nuys,0,0,Fiber Optic,34.178483,-118.43179099999999,1,86.45,0,6,None,40376,1,0,1,1,43,1,0.0,906.44,0.0,3574.5,0,1,91401
1875,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),114.1,8086.4,0,64,3,23.27,4965,0,Fallbrook,1,1,DSL,33.362575,-117.299644,1,114.1,0,6,None,42239,1,0,1,1,72,1,0.0,1675.44,0.0,8086.4,0,1,92028
1876,1,0,1,0,47,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),95.2,4563,0,21,85,20.93,4977,0,Sherman Oaks,0,1,DSL,34.147149,-118.463365,1,95.2,0,1,None,22085,0,0,1,1,47,1,3879.0,983.71,0.0,4563.0,1,0,91403
1877,1,0,0,0,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),88.55,6362.35,0,61,27,46.1,6468,0,Van Nuys,1,1,Cable,34.202494,-118.448048,0,88.55,0,0,None,51348,1,0,0,1,72,1,0.0,3319.2000000000007,0.0,6362.35,0,1,91405
1878,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.75,67.1,0,23,0,16.39,2406,0,Van Nuys,0,1,NA,34.195685,-118.490752,0,20.75,0,0,Offer E,50047,0,0,0,0,3,0,0.0,49.17,0.0,67.1,1,0,91406
1879,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.05,70.05,1,38,22,27.89,2699,1,Van Nuys,0,1,Fiber Optic,34.178470000000004,-118.45947199999999,0,72.852,0,0,None,23646,0,0,0,0,1,4,0.0,27.89,0.0,70.05,0,1,91411
1880,1,0,0,0,2,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.0,165.45,1,61,33,43.47,4546,1,Sherman Oaks,0,1,Cable,34.146957,-118.432138,0,89.44,0,0,Offer E,29387,0,2,0,1,2,3,0.0,86.94,0.0,165.45,0,1,91423
1881,1,0,0,0,26,0,No phone service,DSL,1,1,0,1,Month-to-month,1,Bank transfer (automatic),44.65,1156.55,0,39,6,0.0,4512,0,Encino,0,1,Cable,34.152875,-118.486056,0,44.65,0,0,None,13129,0,2,0,1,26,1,69.0,0.0,0.0,1156.55,0,0,91436
1882,1,0,1,1,29,1,0,DSL,1,0,0,1,Month-to-month,1,Mailed check,60.2,1834.15,0,28,73,1.41,5517,0,Burbank,0,1,DSL,34.188339,-118.30094199999999,1,60.2,3,9,None,18112,0,0,1,1,29,2,0.0,40.89,0.0,1834.15,1,1,91501
1883,0,1,1,0,35,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Bank transfer (automatic),100.5,3653.35,1,65,24,15.98,4745,1,Burbank,0,0,Fiber Optic,34.177267,-118.31003,1,104.52,0,1,None,11517,1,2,1,0,35,6,877.0,559.3000000000002,0.0,3653.35,0,0,91502
1884,1,0,0,0,27,1,0,DSL,1,1,0,0,One year,0,Bank transfer (automatic),55.45,1477.65,0,50,21,20.29,3616,0,Burbank,0,1,Cable,34.213049,-118.317651,0,55.45,0,0,None,25882,0,0,0,0,27,1,0.0,547.8299999999998,0.0,1477.65,0,1,91504
1885,1,0,1,1,24,1,0,DSL,1,1,0,1,Month-to-month,1,Credit card (automatic),70.3,1706.45,0,30,26,44.57,3359,0,Burbank,0,1,Fiber Optic,34.174215000000004,-118.345928,1,70.3,2,6,None,29245,1,1,1,1,24,2,0.0,1069.68,0.0,1706.45,0,1,91505
1886,1,0,1,1,67,1,0,DSL,1,0,0,0,Two year,1,Bank transfer (automatic),60.4,3953.7,0,60,13,21.17,5356,0,Burbank,1,1,Cable,34.169706,-118.323548,1,60.4,0,1,None,18539,1,0,1,0,67,2,51.4,1418.39,0.0,3953.7,0,1,91506
1887,0,0,0,0,16,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,72.65,1194.3,1,35,19,46.99,2850,1,North Hollywood,0,0,DSL,34.1692,-118.372498,0,75.55600000000003,0,0,Offer D,36625,0,2,0,0,16,6,0.0,751.84,0.0,1194.3,0,1,91601
1888,0,0,0,0,23,1,0,DSL,0,1,0,0,One year,0,Bank transfer (automatic),55.8,1327.85,0,55,8,9.04,2499,0,North Hollywood,1,0,Fiber Optic,34.15136,-118.36478600000001,0,55.8,0,0,Offer D,16996,0,0,0,0,23,0,106.0,207.92,0.0,1327.85,0,0,91602
1889,1,0,0,0,14,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Mailed check,31.1,419.7,0,63,12,0.0,3448,0,Studio City,0,1,Fiber Optic,34.139082,-118.39275,0,31.1,0,0,Offer D,26157,0,0,0,0,14,2,0.0,0.0,0.0,419.7,0,1,91604
1890,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,21.0,21,1,30,0,16.66,3753,1,North Hollywood,0,0,NA,34.207295,-118.40002199999999,1,21.0,0,1,Offer E,57146,0,0,1,0,1,4,0.0,16.66,0.0,21.0,0,0,91605
1891,0,1,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.1,45.1,1,80,15,15.24,2740,1,North Hollywood,0,0,DSL,34.187599,-118.387125,0,46.903999999999996,0,0,Offer E,45358,0,2,0,0,1,5,0.0,15.24,0.0,45.1,0,1,91606
1892,1,1,0,0,4,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Credit card (automatic),50.95,207.35,0,72,10,0.0,2104,0,Valley Village,0,1,Fiber Optic,34.165783000000005,-118.399795,0,50.95,0,0,None,27453,0,1,0,0,4,2,2.07,0.0,0.0,207.35,0,1,91607
1893,1,0,0,1,16,1,1,DSL,1,1,0,1,Month-to-month,1,Electronic check,69.1,1083.7,0,46,18,13.99,5172,0,Rancho Cucamonga,0,1,Fiber Optic,34.132275,-117.611478,0,69.1,2,0,Offer D,39064,0,0,0,1,16,1,19.51,223.84,0.0,1083.7,0,1,91701
1894,0,0,1,0,46,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,43.95,2007.85,0,47,8,0.0,4818,0,Azusa,0,0,DSL,34.174493,-117.87068000000001,1,43.95,0,1,None,57775,0,0,1,1,46,0,161.0,0.0,0.0,2007.85,0,0,91702
1895,1,0,0,1,68,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),86.5,5882.75,0,62,29,11.5,4280,0,Baldwin Park,0,1,Fiber Optic,34.098275,-117.967399,0,86.5,0,0,None,76890,1,0,0,1,68,1,0.0,782.0,0.0,5882.75,0,1,91706
1896,1,0,0,0,38,1,1,DSL,1,1,0,0,Month-to-month,0,Electronic check,69.95,2657.55,0,51,22,28.0,5858,0,Chino Hills,1,1,Cable,33.942895,-117.72564399999999,0,69.95,0,0,None,66754,1,0,0,0,38,0,585.0,1064.0,0.0,2657.55,0,0,91709
1897,1,1,1,0,30,1,0,DSL,0,1,0,0,Month-to-month,1,Bank transfer (automatic),50.4,1527.5,1,71,32,4.65,4795,1,Chino,0,1,Fiber Optic,33.990646000000005,-117.663025,1,52.416000000000004,0,1,None,75319,0,0,1,0,30,1,489.0,139.5,0.0,1527.5,0,0,91710
1898,0,1,0,0,5,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,78.95,378.4,1,70,22,12.27,4054,1,Claremont,0,0,Fiber Optic,34.127621000000005,-117.717863,0,82.10799999999999,0,0,Offer E,34716,0,0,0,0,5,5,83.0,61.35,0.0,378.4,0,0,91711
1899,1,0,0,0,17,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),90.95,1612.2,0,49,21,34.98,5687,0,Covina,1,1,DSL,34.097345000000004,-117.90673600000001,0,90.95,0,0,Offer D,33817,0,0,0,1,17,0,339.0,594.66,0.0,1612.2,0,0,91722
1900,1,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.9,76.65,0,25,0,24.57,2347,0,Covina,0,1,NA,34.084747,-117.886844,1,19.9,1,1,Offer E,17554,0,0,1,0,4,0,0.0,98.28,0.0,76.65,1,0,91723
1901,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,20.15,260.7,0,35,0,26.67,4628,0,Covina,0,0,NA,34.081109999999995,-117.853935,0,20.15,0,0,Offer D,25068,0,0,0,0,12,0,0.0,320.04,0.0,260.7,0,0,91724
1902,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),90.6,6441.85,0,57,11,34.97,4528,0,Rancho Cucamonga,1,1,DSL,34.100970000000004,-117.57882,1,90.6,0,1,None,51970,1,0,1,1,72,0,709.0,2517.84,0.0,6441.85,0,0,91730
1903,1,0,0,0,3,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,92.0,266.8,0,58,9,15.6,4345,0,El Monte,0,1,DSL,34.079934,-118.046695,0,92.0,0,0,Offer E,30211,0,0,0,1,3,1,24.0,46.8,0.0,266.8,0,0,91731
1904,1,0,0,0,56,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,94.45,5124.6,1,21,56,25.41,4830,1,El Monte,0,1,Fiber Optic,34.074492,-118.01462,0,98.228,0,0,None,62660,1,0,0,1,56,2,2870.0,1422.96,0.0,5124.6,1,0,91732
1905,0,0,0,0,41,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,24.85,962.25,0,38,0,32.66,3089,0,South El Monte,0,0,NA,34.04622,-118.053753,0,24.85,0,0,None,45645,0,0,0,0,41,0,0.0,1339.06,0.0,962.25,0,0,91733
1906,1,0,0,0,40,0,No phone service,DSL,0,1,0,0,One year,0,Credit card (automatic),36.0,1382.9,0,55,12,0.0,5323,0,Rancho Cucamonga,0,1,DSL,34.245289,-117.642503,0,36.0,0,0,None,23079,1,0,0,0,40,2,166.0,0.0,0.0,1382.9,0,0,91737
1907,0,0,0,0,7,1,0,DSL,1,1,1,1,Month-to-month,1,Electronic check,78.5,571.05,0,44,13,3.34,3601,0,Rancho Cucamonga,0,0,Fiber Optic,34.133809,-117.523724,0,78.5,0,0,Offer E,12937,1,1,0,1,7,1,74.0,23.38,0.0,571.05,0,0,91739
1908,1,0,0,0,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.95,1399.35,0,24,0,7.18,4328,0,Glendora,0,1,NA,34.119363,-117.85505900000001,0,19.95,0,0,None,25135,0,0,0,0,69,2,0.0,495.42,0.0,1399.35,1,0,91740
1909,1,0,1,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.65,150,0,64,0,21.09,2874,0,Glendora,0,1,NA,34.14649,-117.84981499999999,1,20.65,0,1,None,24973,0,0,1,0,7,1,0.0,147.63,0.0,150.0,0,0,91741
1910,0,0,1,1,5,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,30.5,167.2,0,22,59,0.0,5973,0,La Puente,0,0,Fiber Optic,34.031441,-117.93643600000001,1,30.5,1,1,None,84965,0,0,1,0,5,0,99.0,0.0,0.0,167.2,1,0,91744
1911,0,0,1,1,72,1,1,Fiber optic,1,1,1,0,Two year,0,Credit card (automatic),106.1,7657.4,0,57,14,6.41,5146,0,Hacienda Heights,1,0,DSL,33.998471,-117.973758,1,106.1,1,1,None,53686,1,0,1,0,72,3,1072.0,461.52,0.0,7657.4,0,0,91745
1912,1,0,1,1,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.5,865.05,0,64,0,27.4,3093,0,La Puente,0,1,NA,34.038983,-117.991372,1,20.5,0,1,None,30802,0,0,1,0,44,0,0.0,1205.6,0.0,865.05,0,0,91746
1913,0,0,0,0,65,1,1,Fiber optic,0,1,1,0,One year,1,Electronic check,95.5,6153.85,0,59,6,27.68,6153,0,Rowland Heights,1,0,Fiber Optic,33.976753,-117.89736699999999,0,95.5,0,0,None,46342,0,0,0,0,65,1,369.0,1799.2,0.0,6153.85,0,0,91748
1914,0,0,0,0,3,1,1,DSL,0,0,1,0,Month-to-month,0,Electronic check,64.6,174.2,0,20,48,40.99,5277,0,La Verne,0,0,Fiber Optic,34.144703,-117.770299,0,64.6,0,0,None,35530,1,0,0,0,3,0,0.0,122.97,0.0,174.2,1,1,91750
1915,1,0,0,0,24,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),51.1,1269.6,0,45,2,2.33,2515,0,Mira Loma,0,1,Fiber Optic,33.999992,-117.535395,0,51.1,0,0,None,18980,1,0,0,0,24,0,25.0,55.92,0.0,1269.6,0,0,91752
1916,0,0,0,0,44,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),84.8,3862.55,1,54,7,40.17,3997,1,Monterey Park,1,0,Fiber Optic,34.050321999999994,-118.14703700000001,0,88.19200000000001,0,0,None,33280,0,1,0,0,44,1,0.0,1767.48,0.0,3862.55,0,1,91754
1917,0,1,1,0,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.1,6352.4,0,70,13,24.44,4627,0,Monterey Park,1,0,Cable,34.049172,-118.115022,1,89.1,0,1,None,26933,1,0,1,0,72,1,0.0,1759.68,0.0,6352.4,0,1,91755
1918,1,0,0,0,24,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,54.95,1348.5,0,28,69,30.07,3407,0,Mt Baldy,0,1,DSL,34.231318,-117.66203200000001,0,54.95,0,0,None,47,1,0,0,0,24,2,0.0,721.6800000000002,0.0,1348.5,1,1,91759
1919,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.9,50.9,1,50,12,6.95,5111,1,Ontario,1,1,Fiber Optic,34.035602000000004,-117.591528,0,52.93600000000001,0,0,Offer E,56280,0,0,0,0,1,1,0.0,6.95,0.0,50.9,0,0,91761
1920,1,0,1,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.45,471.55,0,43,0,20.78,3727,0,Ontario,0,1,NA,34.057256,-117.667677,1,20.45,0,1,Offer D,54254,0,0,1,0,22,0,0.0,457.16,0.0,471.55,0,0,91762
1921,1,0,1,1,70,1,1,DSL,0,1,1,1,Two year,1,Credit card (automatic),85.95,5931.75,0,33,24,30.06,6354,0,Montclair,1,1,Fiber Optic,34.072121,-117.698319,1,85.95,0,10,None,34447,1,0,1,1,70,1,1424.0,2104.2,0.0,5931.75,0,0,91763
1922,1,0,1,1,25,1,1,DSL,0,0,1,0,Month-to-month,0,Electronic check,60.35,1404.65,0,55,76,25.87,3192,0,Ontario,0,1,Cable,34.074087,-117.60561799999999,1,60.35,3,1,None,49474,0,0,1,0,25,0,0.0,646.75,0.0,1404.65,0,1,91764
1923,1,0,1,1,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.8,726.1,0,24,0,8.21,2745,0,Diamond Bar,0,1,NA,33.992416,-117.807874,1,19.8,3,0,None,46532,0,1,0,0,37,4,0.0,303.7700000000001,0.0,726.1,1,0,91765
1924,0,1,1,1,22,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Bank transfer (automatic),85.35,1961.6,0,71,27,40.19,2656,0,Pomona,0,0,Fiber Optic,34.042286,-117.756106,1,85.35,1,7,Offer D,69974,0,0,1,0,22,1,530.0,884.18,0.0,1961.6,0,0,91766
1925,0,0,1,1,59,1,1,DSL,0,0,1,0,Two year,1,Bank transfer (automatic),72.1,4194.85,0,39,24,24.81,6225,0,Pomona,1,0,Fiber Optic,34.083086,-117.737997,1,72.1,0,9,None,46626,1,0,1,0,59,1,1007.0,1463.79,0.0,4194.85,0,0,91767
1926,1,0,1,1,49,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.8,4872.45,1,27,80,46.94,6088,1,Pomona,1,1,Cable,34.067932,-117.785168,1,103.792,0,1,None,36057,0,0,1,1,49,3,3898.0,2300.06,0.0,4872.45,1,0,91768
1927,1,0,1,1,47,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),107.35,5118.95,1,43,8,37.74,3620,1,Rosemead,1,1,Cable,34.065108,-118.08279099999999,1,111.644,0,1,None,61623,1,1,1,1,47,2,40.95,1773.7800000000002,0.0,5118.95,0,1,91770
1928,0,0,1,1,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.55,658.95,1,45,0,30.07,2687,1,San Dimas,0,0,NA,34.102119,-117.815532,1,19.55,0,1,None,33878,0,2,1,0,31,1,0.0,932.17,0.0,658.95,0,0,91773
1929,1,0,1,1,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,81.05,81.05,0,19,85,36.32,4396,0,San Gabriel,0,1,Cable,34.114771999999995,-118.089431,1,81.05,3,1,None,23444,0,0,1,1,1,0,0.0,36.32,0.0,81.05,1,0,91775
1930,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.5,76.95,0,28,0,37.01,5296,0,San Gabriel,0,1,NA,34.089927,-118.09564499999999,0,20.5,0,0,None,38041,0,0,0,0,3,0,0.0,111.03,0.0,76.95,1,0,91776
1931,0,0,1,0,53,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),111.8,5809.75,0,29,69,41.82,5713,0,Temple City,1,0,Fiber Optic,34.101608,-118.055848,1,111.8,0,3,None,32718,1,0,1,1,53,0,0.0,2216.46,0.0,5809.75,1,1,91780
1932,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.2,20.2,0,27,0,42.15,3586,0,Upland,0,1,NA,34.141146,-117.65558300000001,0,20.2,0,0,None,23331,0,0,0,0,1,1,0.0,42.15,0.0,20.2,1,0,91784
1933,1,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.7,415.9,0,59,0,30.13,2860,0,Upland,0,1,NA,34.105493,-117.66093400000001,0,19.7,0,0,Offer D,48827,0,0,0,0,20,4,0.0,602.6,0.0,415.9,0,0,91786
1934,0,0,0,0,3,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,79.1,246.5,1,60,2,32.43,5339,1,Walnut,0,0,Fiber Optic,34.018353999999995,-117.85491999999999,0,82.264,0,0,Offer E,45118,0,0,0,0,3,3,5.0,97.29,0.0,246.5,0,0,91789
1935,0,0,0,0,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.85,996.95,0,61,0,29.87,5089,0,West Covina,0,0,NA,34.066964,-117.93700700000001,0,19.85,0,0,Offer B,44099,0,0,0,0,51,1,0.0,1523.37,0.0,996.95,0,0,91790
1936,0,0,1,0,51,1,0,DSL,1,1,0,0,One year,1,Bank transfer (automatic),60.5,3145.15,0,56,12,47.18,4207,0,West Covina,0,0,Cable,34.061634000000005,-117.893169,1,60.5,0,4,Offer B,30458,1,0,1,0,51,1,37.74,2406.18,0.0,3145.15,0,1,91791
1937,0,0,1,1,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.55,265.3,0,21,0,42.23,2816,0,West Covina,0,0,NA,34.024405,-117.89872199999999,1,19.55,3,1,None,31622,0,0,1,0,13,2,0.0,548.99,0.0,265.3,1,0,91792
1938,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.9,20.9,0,28,0,10.21,3901,0,Alhambra,0,0,NA,34.090925,-118.12816399999998,0,20.9,0,0,None,54382,0,0,0,0,1,0,0.0,10.21,0.0,20.9,1,0,91801
1939,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,21.05,21.05,0,53,0,10.14,3389,0,Alhambra,0,1,NA,34.074736,-118.145959,0,21.05,1,0,None,30635,0,0,0,0,1,2,0.0,10.14,0.0,21.05,0,0,91803
1940,1,0,0,0,63,1,1,DSL,1,1,0,0,One year,0,Electronic check,71.5,4576.3,0,46,11,18.05,5342,0,Alpine,1,1,Cable,32.827184,-116.70372900000001,0,71.5,0,0,Offer B,16486,1,0,0,0,63,0,50.34,1137.15,0.0,4576.3,0,1,91901
1941,1,0,0,0,3,1,0,DSL,0,0,0,1,Month-to-month,0,Mailed check,54.65,189.1,0,64,30,33.53,2168,0,Bonita,0,1,Fiber Optic,32.671170000000004,-117.00232,0,54.65,0,0,None,17389,0,0,0,1,3,3,57.0,100.59,0.0,189.1,0,0,91902
1942,1,0,0,0,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.2,908.15,0,49,0,30.99,2776,0,Boulevard,0,1,NA,32.677096999999996,-116.30499099999999,0,19.2,0,0,Offer B,1509,0,0,0,0,46,0,0.0,1425.54,0.0,908.15,0,0,91905
1943,1,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),49.8,49.8,0,31,11,3.97,4796,0,Campo,0,1,Fiber Optic,32.673483000000004,-116.47286299999999,0,49.8,0,0,None,3133,0,0,0,0,1,1,0.0,3.97,0.0,49.8,0,1,91906
1944,1,0,0,1,8,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,25.5,215.2,1,40,18,0.0,5578,1,San Diego,0,1,Fiber Optic,32.825086,-117.199424,0,26.52,0,0,None,51213,0,0,0,0,8,5,39.0,0.0,0.0,215.2,0,0,92117
1945,0,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.5,1500.95,0,60,0,11.13,4941,0,Chula Vista,0,0,NA,32.607964,-117.059459,1,20.5,1,8,None,71126,0,0,1,0,71,0,0.0,790.23,0.0,1500.95,0,0,91911
1946,1,0,1,1,55,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),90.4,5099.15,0,38,56,22.56,4603,0,Chula Vista,1,1,Fiber Optic,32.64164,-116.985026,1,90.4,3,10,Offer B,12884,0,0,1,0,55,2,0.0,1240.8,0.0,5099.15,0,1,91913
1947,0,0,0,0,70,1,1,Fiber optic,0,1,0,0,One year,1,Bank transfer (automatic),90.25,6385.95,0,38,3,13.4,5327,0,Chula Vista,1,0,Fiber Optic,32.688506,-116.93863200000001,0,90.25,0,0,None,2606,1,0,0,0,70,0,19.16,938.0,0.0,6385.95,0,1,91914
1948,0,0,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,80.75,159.45,1,41,7,5.11,2176,1,San Diego,0,0,Cable,32.825086,-117.199424,0,83.98,0,0,None,51213,0,0,0,1,2,0,11.0,10.22,0.0,159.45,0,0,92117
1949,1,0,1,1,67,1,1,Fiber optic,1,0,1,1,Two year,0,Bank transfer (automatic),104.6,6885.75,0,32,57,11.31,4743,0,Descanso,0,1,DSL,32.912664,-116.63538700000001,1,104.6,3,10,None,1587,1,0,1,1,67,1,3925.0,757.77,0.0,6885.75,0,0,91916
1950,1,0,1,0,65,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),91.85,5940.85,1,29,80,36.75,5530,1,San Diego,0,1,Cable,32.825086,-117.199424,1,95.524,0,0,None,51213,0,2,0,1,65,5,4753.0,2388.75,0.0,5940.85,1,0,92117
1951,1,0,1,0,14,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),50.2,668.85,0,27,59,4.05,4253,0,Guatay,1,1,Fiber Optic,32.857946000000005,-116.561917,1,50.2,0,6,None,796,0,0,1,0,14,0,395.0,56.7,0.0,668.85,1,0,91931
1952,0,0,1,1,20,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),95.5,1916.2,0,28,48,38.71,3186,0,Imperial Beach,1,0,Cable,32.579134,-117.119009,1,95.5,2,5,None,26662,1,0,1,1,20,0,920.0,774.2,0.0,1916.2,1,0,91932
1953,1,0,0,1,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,75.35,75.35,1,41,23,32.82,5284,1,San Diego,0,1,Fiber Optic,32.825086,-117.199424,0,78.36399999999998,0,0,None,51213,0,0,0,0,1,5,0.0,32.82,0.0,75.35,0,0,92117
1954,1,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.45,75.45,1,55,16,11.58,5518,1,San Diego,0,1,Cable,32.825086,-117.199424,0,78.468,0,0,None,51213,0,2,0,0,1,5,0.0,11.58,0.0,75.45,0,0,92117
1955,0,0,1,1,49,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.4,4613.95,0,56,53,8.18,6136,0,La Mesa,0,0,Cable,32.759327,-116.99726000000001,1,95.4,6,6,Offer B,44652,0,1,1,1,49,2,2445.0,400.82,0.0,4613.95,0,0,91941
1956,0,0,0,0,72,1,1,Fiber optic,1,1,1,0,Two year,1,Bank transfer (automatic),101.3,7261.25,0,32,16,2.25,5513,0,La Mesa,1,0,Cable,32.782501,-117.01611000000001,0,101.3,0,0,Offer A,24005,0,0,0,0,72,0,0.0,162.0,0.0,7261.25,0,1,91942
1957,0,0,1,0,46,1,1,DSL,1,0,0,0,Month-to-month,0,Electronic check,53.1,2459.8,0,25,82,44.74,3358,0,Lemon Grove,0,0,Fiber Optic,32.733564,-117.03371299999999,1,53.1,0,1,Offer B,24961,0,0,1,1,46,0,201.7,2058.04,0.0,2459.8,1,1,91945
1958,1,0,0,0,24,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),84.85,2048.8,0,57,14,13.13,2941,0,Mount Laguna,1,1,Fiber Optic,32.830852,-116.444601,0,84.85,0,0,Offer C,81,0,0,0,0,24,0,28.68,315.12,0.0,2048.8,0,1,91948
1959,0,0,1,1,5,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,34.25,163.55,0,52,19,0.0,5100,0,National City,0,0,DSL,32.67102,-117.095235,1,34.25,2,9,None,62355,1,0,1,0,5,0,0.0,0.0,0.0,163.55,0,1,91950
1960,0,0,1,1,33,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Credit card (automatic),88.6,2888.7,0,21,73,11.01,3648,0,Pine Valley,1,0,Fiber Optic,32.800671,-116.48336299999998,1,88.6,1,6,Offer C,1604,1,0,1,1,33,1,2109.0,363.33,0.0,2888.7,1,0,91962
1961,0,0,0,0,42,1,1,DSL,1,1,0,0,One year,1,Bank transfer (automatic),60.15,2421.6,0,23,41,29.44,5988,0,Potrero,0,0,Fiber Optic,32.619465000000005,-116.59360500000001,0,60.15,0,0,Offer B,905,0,0,0,1,42,0,993.0,1236.48,0.0,2421.6,1,0,91963
1962,1,0,0,0,23,1,0,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),99.95,2292.75,0,21,30,41.94,3515,0,Spring Valley,1,1,DSL,32.726627,-116.99460800000001,0,99.95,0,0,None,56100,0,0,0,1,23,1,688.0,964.62,0.0,2292.75,1,0,91977
1963,1,0,0,0,8,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),70.7,553.4,0,26,59,41.93,4946,0,Spring Valley,0,1,DSL,32.730264,-116.95096299999999,0,70.7,0,0,Offer E,7863,0,0,0,1,8,3,0.0,335.44,0.0,553.4,1,1,91978
1964,1,0,0,0,66,1,0,DSL,1,1,0,0,One year,1,Mailed check,54.8,3465.7,0,32,30,11.56,4621,0,Tecate,0,1,DSL,32.587557000000004,-116.636816,0,54.8,0,0,Offer A,91,0,0,0,0,66,0,0.0,762.96,0.0,3465.7,0,1,91980
1965,1,0,0,0,24,1,0,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),49.55,1210.4,1,35,31,14.39,5005,1,San Diego,0,1,Cable,32.825086,-117.199424,0,51.532,0,0,None,51213,0,1,0,0,24,1,375.0,345.36,0.0,1210.4,0,0,92117
1966,1,1,0,0,24,1,1,DSL,0,1,0,0,Month-to-month,0,Credit card (automatic),54.8,1291.3,0,74,27,8.66,4330,0,Borrego Springs,0,1,Fiber Optic,33.200369,-116.19231299999998,0,54.8,0,0,None,2863,0,0,0,0,24,0,349.0,207.84,0.0,1291.3,0,0,92004
1967,1,0,0,0,69,1,1,DSL,1,1,0,1,One year,1,Credit card (automatic),78.6,5356.45,1,51,10,29.38,6230,1,San Diego,1,1,Fiber Optic,32.825086,-117.199424,0,81.744,0,0,Offer A,51213,1,0,0,1,69,1,536.0,2027.22,0.0,5356.45,0,0,92117
1968,0,0,0,0,53,1,0,Fiber optic,0,1,1,1,One year,1,Mailed check,100.3,5200.8,0,22,73,8.33,5377,0,Carlsbad,1,0,DSL,33.148115999999995,-117.30604299999999,0,100.3,0,0,Offer B,35582,0,0,0,1,53,2,3797.0,441.49,0.0,5200.8,1,0,92008
1969,0,0,0,0,60,0,No phone service,DSL,1,0,1,1,Two year,0,Electronic check,53.6,3237.05,0,61,4,0.0,4173,0,Carlsbad,1,0,DSL,33.098017999999996,-117.25820300000001,0,53.6,0,0,None,43161,0,1,0,1,60,1,0.0,0.0,0.0,3237.05,0,1,92009
1970,0,0,1,0,7,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,81.1,576.65,1,35,30,11.58,3238,1,San Diego,0,0,Cable,32.825086,-117.199424,1,84.344,0,1,None,51213,0,0,1,0,7,3,173.0,81.06,0.0,576.65,0,0,92117
1971,0,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),19.35,433.75,0,32,0,10.9,5811,0,El Cajon,0,0,NA,32.785165,-116.862648,0,19.35,0,0,None,40995,0,2,0,0,20,1,0.0,218.0,0.0,433.75,0,0,92019
1972,0,0,1,1,23,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,85.6,1868.4,0,25,71,9.84,3513,0,El Cajon,0,0,DSL,32.79697,-116.969082,1,85.6,1,10,None,55277,0,0,1,1,23,1,0.0,226.32,0.0,1868.4,1,1,92020
1973,1,0,1,1,72,1,0,DSL,1,0,1,1,Two year,1,Electronic check,80.8,5728.55,0,23,53,35.07,4689,0,El Cajon,1,1,Fiber Optic,32.832706,-116.873258,1,80.8,0,8,Offer A,61872,1,0,1,1,72,1,303.61,2525.04,0.0,5728.55,1,1,92021
1974,1,0,1,0,11,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.95,825.7,1,39,33,21.58,2044,1,San Diego,0,1,Cable,32.825086,-117.199424,1,77.94800000000002,0,1,Offer D,51213,0,0,1,0,11,1,272.0,237.38,0.0,825.7,0,0,92117
1975,1,0,0,0,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.6,390.4,0,43,0,16.81,4562,0,Escondido,0,1,NA,33.081478000000004,-117.03381399999999,0,19.6,0,0,None,49281,0,0,0,0,21,0,0.0,353.01,0.0,390.4,0,0,92025
1976,1,1,0,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.55,93.55,1,73,7,30.17,5536,1,San Diego,0,1,DSL,32.825086,-117.199424,0,97.292,0,0,Offer E,51213,0,1,0,0,1,4,0.0,30.17,0.0,93.55,0,0,92117
1977,1,1,0,0,31,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,90.7,2845.15,0,75,24,46.71,3493,0,Escondido,0,1,Fiber Optic,33.141265000000004,-116.967221,0,90.7,0,0,None,48690,0,0,0,0,31,0,683.0,1448.01,0.0,2845.15,0,0,92027
1978,0,0,0,0,57,1,0,DSL,0,1,1,0,Two year,0,Mailed check,69.75,3894.4,0,21,48,36.14,4487,0,Fallbrook,1,0,Fiber Optic,33.362575,-117.299644,0,69.75,0,0,None,42239,1,0,0,1,57,0,1869.0,2059.98,0.0,3894.4,1,0,92028
1979,0,0,1,1,45,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.0,886.4,0,42,0,21.73,5169,0,Escondido,0,0,NA,33.079834000000005,-117.134275,1,20.0,2,9,None,17944,0,0,1,0,45,1,0.0,977.85,0.0,886.4,0,0,92029
1980,1,0,0,0,10,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,95.25,1021.55,0,35,13,26.43,4810,0,Julian,1,1,Fiber Optic,32.980678000000005,-116.262854,0,95.25,0,0,None,3577,0,1,0,1,10,1,133.0,264.3,0.0,1021.55,0,0,92036
1981,0,0,1,0,58,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),102.1,5885.4,1,33,31,3.51,4415,1,San Diego,1,0,Cable,32.825086,-117.199424,1,106.184,0,1,None,51213,1,2,1,1,58,2,1824.0,203.58,0.0,5885.4,0,0,92117
1982,1,0,0,1,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,268.4,0,49,0,40.66,5770,0,Lakeside,0,1,NA,32.909873,-116.906774,0,19.95,5,0,None,42277,0,0,0,0,14,2,0.0,569.24,0.0,268.4,0,0,92040
1983,1,0,1,0,27,1,1,DSL,1,0,1,1,One year,0,Mailed check,80.85,2204.35,0,42,14,11.83,4732,0,Oceanside,0,1,DSL,33.351059,-117.420557,1,80.85,0,3,Offer C,98239,1,0,1,1,27,1,0.0,319.41,0.0,2204.35,0,1,92054
1984,0,0,1,1,14,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),90.9,1259,1,64,10,13.64,5148,1,San Diego,0,0,DSL,32.825086,-117.199424,1,94.53600000000002,0,1,Offer D,51213,0,0,1,1,14,1,126.0,190.96,0.0,1259.0,0,0,92117
1985,0,0,1,1,12,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Mailed check,29.2,309.1,1,46,30,0.0,3747,1,San Diego,0,0,Cable,32.825086,-117.199424,1,30.368000000000002,0,1,None,51213,0,2,1,0,12,4,0.0,0.0,0.0,309.1,0,1,92117
1986,0,0,1,1,69,1,1,Fiber optic,0,1,0,1,Two year,1,Bank transfer (automatic),93.3,6398.05,0,59,24,28.53,5205,0,Pala,0,0,Fiber Optic,33.384345,-117.07261899999999,1,93.3,1,0,Offer A,1831,1,0,0,1,69,2,1536.0,1968.57,0.0,6398.05,0,0,92059
1987,0,0,1,1,25,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),89.15,2257.75,1,36,6,24.64,5853,1,San Diego,1,0,Fiber Optic,32.825086,-117.199424,1,92.716,0,1,None,51213,0,1,1,0,25,1,0.0,616.0,0.0,2257.75,0,1,92117
1988,1,1,1,0,58,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,108.85,6287.25,1,78,21,49.38,4739,1,San Diego,1,1,Fiber Optic,32.825086,-117.199424,1,113.204,0,1,None,51213,0,0,1,0,58,0,1320.0,2864.04,0.0,6287.25,0,0,92117
1989,0,0,1,1,35,0,No phone service,DSL,1,0,1,0,Two year,1,Credit card (automatic),46.35,1662.05,0,59,24,0.0,4577,0,Poway,0,0,DSL,32.984395,-117.01345400000001,1,46.35,0,7,Offer C,47969,1,0,1,0,35,0,39.89,0.0,0.0,1662.05,0,1,92064
1990,0,1,0,0,16,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.75,1350.15,1,76,8,17.51,5136,1,San Diego,0,0,Fiber Optic,32.825086,-117.199424,0,88.14,0,0,None,51213,0,2,0,0,16,8,108.0,280.16,0.0,1350.15,0,0,92117
1991,1,0,1,1,45,1,1,DSL,0,1,1,1,One year,0,Credit card (automatic),78.75,3600.65,0,33,13,39.82,2595,0,Ranchita,1,1,Cable,33.215251,-116.53633,1,78.75,0,3,None,339,0,0,1,1,45,0,468.0,1791.9,0.0,3600.65,0,0,92066
1992,0,0,0,0,17,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,83.55,1329.15,0,60,19,22.61,5564,0,Rancho Santa Fe,0,0,Fiber Optic,33.012751,-117.200617,0,83.55,0,0,None,7615,0,0,0,0,17,1,25.25,384.37,0.0,1329.15,0,1,92067
1993,0,0,1,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.7,45.7,1,37,6,12.8,3187,1,San Diego,0,0,DSL,32.825086,-117.199424,1,47.52800000000001,0,3,None,51213,0,0,1,0,1,2,0.0,12.8,0.0,45.7,0,0,92117
1994,1,0,0,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.6,422.5,0,62,0,20.46,2203,0,Santa Ysabel,0,1,NA,33.174725,-116.743329,0,19.6,0,0,None,1143,0,0,0,0,22,1,0.0,450.12,0.0,422.5,0,0,92070
1995,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.95,69.95,1,73,30,22.5,3208,1,San Diego,0,0,Cable,32.825086,-117.199424,0,72.748,0,0,Offer E,51213,0,0,0,0,1,2,0.0,22.5,0.0,69.95,0,0,92117
1996,1,0,1,1,67,1,0,DSL,1,0,0,1,Two year,0,Mailed check,67.85,4627.65,0,21,58,2.12,4792,0,Solana Beach,1,1,Fiber Optic,33.001813,-117.263628,1,67.85,0,5,Offer A,12173,1,0,1,1,67,1,0.0,142.04000000000005,0.0,4627.65,1,1,92075
1997,0,0,1,1,67,1,1,Fiber optic,0,0,1,1,Two year,1,Bank transfer (automatic),105.65,6717.9,0,45,22,17.79,6383,0,San Marcos,1,0,Fiber Optic,33.119028,-117.166036,1,105.65,3,8,Offer A,6760,1,0,1,1,67,3,1478.0,1191.9299999999996,0.0,6717.9,0,0,92078
1998,0,0,1,0,2,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Electronic check,44.6,97.1,1,23,56,0.0,5482,1,San Diego,0,0,DSL,32.825086,-117.199424,1,46.38399999999999,0,1,None,51213,0,1,1,1,2,2,54.0,0.0,0.0,97.1,1,0,92117
1999,1,0,0,0,23,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.95,1710.45,1,48,14,28.8,5897,1,San Diego,0,1,Fiber Optic,32.825086,-117.199424,0,77.94800000000002,0,0,None,51213,0,0,0,0,23,3,239.0,662.4,0.0,1710.45,0,0,92117
2000,0,1,0,0,9,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),75.5,637.4,0,65,9,24.96,3021,0,Vista,1,0,DSL,33.22784,-117.200024,0,75.5,0,0,None,44692,0,2,0,0,9,3,57.0,224.64,0.0,637.4,0,0,92084
2001,0,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.15,117.95,0,30,0,3.37,5020,0,Warner Springs,0,0,NA,33.323705,-116.626907,0,20.15,0,0,Offer E,1205,0,0,0,0,5,0,0.0,16.85,0.0,117.95,0,0,92086
2002,1,0,0,0,54,0,No phone service,DSL,1,0,1,0,Two year,0,Credit card (automatic),45.2,2460.55,0,47,10,0.0,5435,0,Rancho Santa Fe,0,1,DSL,32.993559999999995,-117.207121,0,45.2,0,0,None,1072,1,0,0,0,54,1,246.0,0.0,0.0,2460.55,0,0,92091
2003,0,0,0,0,57,1,0,Fiber optic,0,0,1,1,Two year,1,Electronic check,95.25,5464.65,1,39,16,17.55,5789,1,San Diego,1,0,DSL,32.825086,-117.199424,0,99.06,0,0,None,51213,0,1,0,1,57,4,874.0,1000.35,0.0,5464.65,0,0,92117
2004,1,0,0,0,24,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,89.85,2165.05,1,23,64,27.97,2050,1,San Diego,1,1,Cable,32.825086,-117.199424,0,93.444,0,0,None,51213,0,0,0,1,24,0,1386.0,671.28,0.0,2165.05,1,0,92117
2005,0,0,1,1,49,1,1,Fiber optic,0,1,1,1,One year,0,Mailed check,100.45,4941.8,1,35,21,26.37,4235,1,San Diego,0,0,DSL,32.825086,-117.199424,1,104.46799999999999,0,1,None,51213,0,0,1,1,49,1,1038.0,1292.13,0.0,4941.8,0,0,92117
2006,1,0,0,0,5,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,47.15,223.15,1,25,94,22.01,2857,1,San Diego,0,1,DSL,32.825086,-117.199424,0,49.036,0,0,None,51213,0,0,0,1,5,5,210.0,110.05,0.0,223.15,1,0,92117
2007,1,0,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.2,181.1,1,58,11,26.47,2384,1,San Diego,0,1,Cable,32.825086,-117.199424,0,83.40799999999999,0,0,None,51213,0,0,0,1,2,5,1.99,52.94,0.0,181.1,0,1,92117
2008,0,0,0,1,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,87.1,341.45,1,33,3,32.46,5587,1,San Diego,1,0,DSL,32.825086,-117.199424,0,90.584,0,0,None,51213,1,2,0,0,4,1,10.0,129.84,0.0,341.45,0,0,92117
2009,1,0,1,1,70,1,1,DSL,1,1,1,0,Two year,1,Bank transfer (automatic),79.25,5731.85,0,56,2,27.97,5085,0,San Diego,1,1,Fiber Optic,32.741852,-117.243453,1,79.25,0,8,Offer A,27959,1,0,1,0,70,2,115.0,1957.9,0.0,5731.85,0,0,92107
2010,1,0,0,0,5,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.9,357.75,1,30,65,46.88,3520,1,San Diego,0,1,DSL,32.825086,-117.199424,0,78.936,0,0,None,51213,0,0,0,0,5,5,233.0,234.4,0.0,357.75,0,0,92117
2011,1,0,1,1,53,1,1,DSL,1,0,1,1,Month-to-month,0,Electronic check,85.7,4616.1,0,51,12,26.84,5957,0,San Diego,1,1,DSL,32.787836,-117.232376,1,85.7,2,5,None,46086,1,2,1,1,53,2,0.0,1422.52,0.0,4616.1,0,1,92109
2012,0,0,1,0,47,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,98.75,4533.7,1,29,56,2.87,4622,1,San Diego,1,0,Cable,32.825086,-117.199424,1,102.7,0,1,None,51213,0,0,1,1,47,4,0.0,134.89,0.0,4533.7,1,1,92117
2013,0,0,0,1,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.1,589.25,0,63,0,33.71,3086,0,San Diego,0,0,NA,32.805518,-117.16905200000001,0,20.1,0,0,Offer C,46828,0,0,0,0,31,2,0.0,1045.01,0.0,589.25,0,0,92111
2014,1,0,1,1,13,1,0,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),61.8,750.1,0,56,56,28.15,4749,0,San Diego,1,1,DSL,32.697098,-117.11658700000001,1,61.8,3,8,None,47431,1,1,1,0,13,2,420.0,365.95,0.0,750.1,0,0,92113
2015,0,0,1,1,28,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,49.9,1410.25,0,33,30,41.41,5250,0,San Diego,0,0,Fiber Optic,32.707892,-117.05512,1,49.9,1,6,Offer C,66838,0,0,1,0,28,1,423.0,1159.48,0.0,1410.25,0,0,92114
2016,0,0,0,0,10,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,86.45,830.85,1,57,22,17.65,5699,1,San Diego,0,0,Fiber Optic,32.825086,-117.199424,0,89.90799999999999,0,0,None,51213,0,0,0,1,10,3,183.0,176.5,0.0,830.85,0,0,92117
2017,1,0,1,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.4,743.5,0,62,0,6.97,3756,0,San Diego,0,1,NA,32.765299,-117.122565,1,20.4,0,8,Offer C,33083,0,1,1,0,38,1,0.0,264.86,0.0,743.5,0,0,92116
2018,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.3,45.3,1,28,65,39.94,3049,1,San Diego,0,0,Cable,32.825086,-117.199424,0,47.111999999999995,0,0,None,51213,0,0,0,1,1,0,0.0,39.94,0.0,45.3,1,0,92117
2019,1,0,1,0,67,1,1,Fiber optic,0,1,1,1,One year,0,Electronic check,104.1,7040.85,1,61,3,8.18,4857,1,Coronado,1,1,Cable,32.68674,-117.18661200000001,1,108.264,0,4,Offer A,24093,0,3,1,1,67,3,0.0,548.06,0.0,7040.85,0,1,92118
2020,1,0,1,0,52,1,0,DSL,1,1,1,1,One year,1,Mailed check,75.4,3865.45,0,28,85,10.4,5211,0,San Diego,0,1,DSL,32.802959,-117.02709499999999,1,75.4,0,9,None,21866,0,0,1,1,52,0,0.0,540.8000000000002,0.0,3865.45,1,1,92119
2021,1,0,1,1,62,1,0,Fiber optic,1,1,1,1,Two year,0,Mailed check,108.15,6825.65,0,42,20,1.76,5298,0,San Diego,1,1,Fiber Optic,32.807867,-117.060993,1,108.15,3,2,None,25569,1,0,1,1,62,0,1365.0,109.12,0.0,6825.65,0,0,92120
2022,0,0,0,0,16,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,86.25,1340.1,0,40,28,22.3,3511,0,San Diego,0,0,DSL,32.898613,-117.202937,0,86.25,0,0,Offer D,4258,0,0,0,1,16,0,0.0,356.8,0.0,1340.1,0,1,92121
2023,0,1,1,0,5,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,81.0,371.65,1,68,12,47.28,4287,1,San Diego,0,0,DSL,32.85723,-117.209774,1,84.24000000000002,0,1,Offer E,34902,0,1,1,0,5,4,0.0,236.4,40.64,371.65,0,1,92122
2024,1,0,0,0,12,1,0,Fiber optic,0,0,1,1,One year,0,Electronic check,95.7,1184,0,57,23,49.0,5527,0,San Diego,1,1,Fiber Optic,32.808814,-117.134694,0,95.7,0,0,Offer D,25232,0,1,0,1,12,2,0.0,588.0,0.0,1184.0,0,1,92123
2025,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),116.85,8477.7,0,63,14,31.83,4055,0,San Diego,1,0,Fiber Optic,32.827238,-117.08928700000001,1,116.85,1,1,Offer A,30206,1,0,1,1,72,0,1187.0,2291.76,0.0,8477.7,0,0,92124
2026,1,1,0,0,71,1,1,Fiber optic,0,1,1,1,One year,0,Bank transfer (automatic),105.75,7382.85,0,80,9,6.1,4921,0,San Diego,0,1,DSL,32.886925,-117.152162,0,105.75,0,0,None,74232,1,0,0,0,71,2,664.0,433.1,0.0,7382.85,0,0,92126
2027,0,0,1,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.15,456.85,0,33,0,32.86,3573,0,San Diego,0,0,NA,33.017518,-117.11845600000001,1,20.15,0,1,Offer C,20046,0,0,1,0,24,2,0.0,788.64,0.0,456.85,0,0,92127
2028,0,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.6,331.6,0,64,0,39.49,2722,0,San Diego,0,0,NA,33.000269,-117.072093,0,19.6,0,0,Offer D,42733,0,0,0,0,15,1,0.0,592.35,0.0,331.6,0,0,92128
2029,1,0,1,0,67,1,0,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),90.6,6056.15,1,31,6,30.75,4394,1,San Diego,0,1,Cable,32.961064,-117.13491699999999,1,94.22399999999999,0,1,Offer A,47224,0,0,1,1,67,1,363.0,2060.25,0.0,6056.15,0,0,92129
2030,1,0,0,1,2,1,1,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),60.95,134.6,0,54,12,14.88,3172,0,San Diego,0,1,Fiber Optic,32.957195,-117.202542,0,60.95,2,0,None,28201,0,0,0,0,2,3,0.0,29.76,0.0,134.6,0,1,92130
2031,0,0,1,1,5,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,25.05,125.5,0,40,53,0.0,2071,0,San Diego,0,0,Fiber Optic,32.89325,-117.08709099999999,1,25.05,3,3,Offer E,29283,0,0,1,0,5,0,0.0,0.0,0.0,125.5,0,1,92131
2032,0,0,1,0,15,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,88.15,1390.6,1,21,84,12.27,2524,1,San Diego,0,0,Cable,32.677716,-117.04766599999999,1,91.67600000000002,0,1,None,36351,0,0,1,1,15,0,0.0,184.05,0.0,1390.6,1,1,92139
2033,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.2,20.2,1,55,0,13.27,4325,1,San Diego,0,1,NA,32.578103000000006,-117.012975,0,20.2,0,0,None,68776,0,0,0,0,1,2,0.0,13.27,0.0,20.2,0,0,92154
2034,1,0,1,1,41,1,0,DSL,1,1,0,0,One year,1,Bank transfer (automatic),60.3,2511.3,0,20,69,2.43,4565,0,San Ysidro,1,1,DSL,32.555828000000005,-117.04007299999999,1,60.3,0,8,None,28488,0,0,1,1,41,0,173.28,99.63,0.0,2511.3,1,1,92173
2035,0,0,0,1,43,1,0,DSL,1,1,0,1,Month-to-month,1,Electronic check,63.95,2737.05,0,26,30,5.6,4205,0,Indio,0,0,DSL,33.713891,-116.237257,0,63.95,1,0,None,56307,0,0,0,1,43,1,821.0,240.8,0.0,2737.05,1,0,92201
2036,1,1,1,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,74.3,74.3,0,76,20,17.84,2968,0,Indio,0,1,DSL,33.752938,-116.23005500000001,1,74.3,0,7,None,2743,0,0,1,0,1,2,0.0,17.84,0.0,74.3,0,0,92203
2037,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.6,70.6,0,73,27,32.61,2576,0,Indian Wells,0,0,Cable,33.537646,-116.29108899999999,0,70.6,0,0,Offer E,3873,0,0,0,0,1,0,0.0,32.61,0.0,70.6,0,1,92210
2038,0,0,1,1,26,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.8,2361.8,1,47,12,15.37,2641,1,Palm Desert,0,0,Cable,33.762759,-116.324817,1,94.432,0,1,None,19702,0,2,1,1,26,6,0.0,399.62,0.0,2361.8,0,1,92211
2039,1,0,0,0,22,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.35,1730.35,1,48,19,19.19,4718,1,Banning,0,1,Cable,33.936298,-116.849577,0,82.524,0,0,None,25859,0,2,0,0,22,5,329.0,422.18,0.0,1730.35,0,0,92220
2040,1,0,1,0,71,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),90.55,6404,0,30,30,28.58,5007,0,Beaumont,1,1,DSL,33.946982,-116.977672,1,90.55,0,2,Offer A,17721,1,0,1,1,71,1,1921.0,2029.18,0.0,6404.0,0,0,92223
2041,1,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.45,165.35,0,29,0,9.43,2600,0,Blythe,0,1,NA,33.674583,-114.71611999999999,0,19.45,0,0,None,24659,0,0,0,0,7,1,0.0,66.00999999999999,0.0,165.35,1,0,92225
2042,0,1,0,0,28,1,1,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),64.45,1867.6,0,67,23,12.72,3820,0,Brawley,1,0,Cable,33.03933,-115.19185700000001,0,64.45,0,0,None,23394,1,0,0,0,28,1,42.95,356.16,0.0,1867.6,0,1,92227
2043,1,1,0,0,16,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.65,1043.3,0,66,24,22.9,5610,0,Cabazon,0,1,Fiber Optic,33.929812,-116.76058,0,69.65,0,0,Offer D,2355,0,0,0,0,16,2,0.0,366.4,0.0,1043.3,0,1,92230
2044,1,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.5,128.6,0,48,0,30.58,4271,0,Calexico,0,1,NA,32.690653999999995,-115.431225,0,19.5,0,0,Offer E,27804,0,0,0,0,7,0,0.0,214.06,0.0,128.6,0,0,92231
2045,0,0,0,0,69,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),110.5,7455.45,0,30,42,23.92,4803,0,Calipatria,1,0,Cable,33.143826000000004,-115.49748500000001,0,110.5,0,0,Offer A,7857,1,0,0,1,69,1,3131.0,1650.48,0.0,7455.45,0,0,92233
2046,0,0,0,1,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,24.7,24.7,0,29,48,0.0,3065,0,Cathedral City,0,0,Fiber Optic,33.829583,-116.474131,0,24.7,1,0,Offer E,43141,0,1,0,0,1,2,0.0,0.0,0.0,24.7,1,1,92234
2047,1,0,0,0,3,1,0,DSL,1,0,1,1,Month-to-month,1,Electronic check,77.4,206.15,0,36,6,44.42,5528,0,Coachella,1,1,Fiber Optic,33.680031,-116.171678,0,77.4,0,0,Offer E,23170,0,0,0,1,3,0,0.0,133.26,0.0,206.15,0,1,92236
2048,1,1,0,0,21,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),96.8,2030.3,1,79,8,42.27,4317,1,Desert Center,1,1,Cable,33.889604999999996,-115.25700900000001,0,100.67200000000001,0,0,None,964,0,1,0,0,21,1,162.0,887.6700000000002,10.2,2030.3,0,0,92239
2049,0,0,1,0,69,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),85.4,5869.4,0,33,29,34.49,5976,0,Desert Hot Springs,1,0,Fiber Optic,33.948558,-116.516976,1,85.4,0,6,Offer A,22796,0,0,1,0,69,0,1702.0,2379.81,0.0,5869.4,0,0,92240
2050,0,0,1,0,71,0,No phone service,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),47.6,3377.8,0,44,16,0.0,4795,0,Desert Hot Springs,1,0,Fiber Optic,33.832799,-116.250973,1,47.6,0,1,Offer A,5529,1,0,1,0,71,1,54.04,0.0,0.0,3377.8,0,1,92241
2051,0,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.4,1346.2,0,19,0,25.18,6408,0,Earp,0,0,NA,34.137741999999996,-114.36514,1,19.4,2,0,Offer A,1564,0,0,0,0,69,0,0.0,1737.42,0.0,1346.2,1,0,92242
2052,0,0,0,0,48,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,103.85,4946.05,0,35,12,10.5,4304,0,El Centro,1,0,Fiber Optic,32.770393,-115.60915,0,103.85,0,0,None,43712,1,0,0,1,48,2,594.0,504.0,0.0,4946.05,0,0,92243
2053,1,0,1,0,47,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),83.35,4065,1,26,65,17.54,2516,1,Heber,1,1,Fiber Optic,32.730583,-115.50108300000001,1,86.684,0,1,Offer B,3535,0,0,1,1,47,0,0.0,824.38,0.0,4065.0,1,1,92249
2054,0,0,0,0,2,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.4,106.55,1,27,57,24.83,5115,1,Fallbrook,0,0,Cable,33.362575,-117.299644,0,51.376000000000005,0,0,None,42239,0,0,0,1,2,0,61.0,49.66,0.0,106.55,1,0,92028
2055,1,0,0,0,45,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Credit card (automatic),108.45,4964.7,0,30,73,5.97,5093,0,Imperial,1,1,Fiber Optic,32.858595,-115.662709,0,108.45,0,0,None,14546,1,0,0,1,45,1,0.0,268.65,0.0,4964.7,0,1,92251
2056,1,0,0,0,51,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),81.0,4085.75,0,54,11,42.93,4121,0,Joshua Tree,0,1,DSL,34.167235999999995,-116.28151100000001,0,81.0,0,0,None,8141,0,0,0,0,51,0,449.0,2189.43,0.0,4085.75,0,0,92252
2057,0,0,1,0,22,1,1,DSL,1,0,1,1,Month-to-month,1,Electronic check,79.2,1742.75,1,27,56,13.11,3410,1,La Quinta,0,0,Cable,33.695532,-116.310571,1,82.36800000000002,0,1,None,23971,1,1,1,1,22,2,976.0,288.42,0.0,1742.75,1,0,92253
2058,1,0,0,0,72,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),86.65,6224.8,0,39,17,11.41,4621,0,Mecca,1,1,DSL,33.543834999999994,-115.99390600000001,0,86.65,0,0,Offer A,8768,1,0,0,1,72,1,0.0,821.52,0.0,6224.8,0,1,92254
2059,1,0,1,1,37,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,92.95,3415.25,0,33,29,38.89,3462,0,Morongo Valley,1,1,DSL,34.097863000000004,-116.59456100000001,1,92.95,1,1,Offer C,3499,0,0,1,0,37,0,0.0,1438.93,0.0,3415.25,0,1,92256
2060,1,0,1,1,71,1,1,DSL,1,1,1,1,Two year,0,Electronic check,90.35,6325.25,0,31,29,18.42,6483,0,Niland,1,1,DSL,33.345825,-115.596574,1,90.35,0,1,Offer A,2753,1,0,1,1,71,3,1834.0,1307.8200000000004,0.0,6325.25,0,0,92257
2061,1,0,1,1,7,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,48.7,340.25,1,61,4,5.13,2984,1,North Palm Springs,1,1,Cable,33.906496000000004,-116.569499,1,50.648,0,1,None,732,0,0,1,0,7,1,14.0,35.91,0.0,340.25,0,0,92258
2062,0,0,0,0,66,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.15,1683.6,0,51,0,20.77,6141,0,Ocotillo,0,0,NA,32.698964000000004,-115.886656,0,25.15,0,0,Offer A,471,0,0,0,0,66,0,0.0,1370.82,0.0,1683.6,0,0,92259
2063,1,0,1,1,51,1,0,DSL,1,0,1,1,One year,1,Bank transfer (automatic),76.4,3966.3,0,59,3,31.66,6385,0,Palm Desert,0,1,DSL,33.694501,-116.41271100000002,1,76.4,0,1,None,29340,1,0,1,1,51,3,11.9,1614.66,0.0,3966.3,0,1,92260
2064,0,0,1,1,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.55,608.5,0,57,0,21.14,5203,0,Palm Springs,0,0,NA,33.839989,-116.65921499999999,1,19.55,0,1,None,24924,0,0,1,0,30,0,0.0,634.2,0.0,608.5,0,0,92262
2065,0,0,0,0,34,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,85.35,2896.6,0,26,76,23.54,3818,0,Palm Springs,0,0,DSL,33.745746000000004,-116.514215,0,85.35,0,0,None,18884,0,0,0,0,34,1,0.0,800.36,0.0,2896.6,1,1,92264
2066,1,0,1,1,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.8,1514.85,0,62,0,35.25,6281,0,Palo Verde,0,1,NA,33.3249,-114.758334,1,24.8,1,1,None,291,0,0,1,0,64,0,0.0,2256.0,0.0,1514.85,0,0,92266
2067,1,1,1,0,65,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),103.15,6792.45,0,65,5,16.65,6441,0,Parker Dam,1,1,Fiber Optic,34.273872,-114.192901,1,103.15,0,1,None,131,0,0,1,1,65,2,0.0,1082.25,0.0,6792.45,0,1,92267
2068,1,0,0,0,47,1,1,Fiber optic,1,1,1,0,Month-to-month,0,Mailed check,100.75,4669.2,0,50,25,47.73,2508,0,Pioneertown,0,1,Fiber Optic,34.201108000000005,-116.593456,0,100.75,0,0,None,354,1,0,0,0,47,1,116.73,2243.31,0.0,4669.2,0,1,92268
2069,0,0,0,0,1,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,95.6,95.6,1,29,30,6.67,4091,1,Rancho Mirage,0,0,Cable,33.763678000000006,-116.429928,0,99.424,0,0,None,12465,0,2,0,1,1,6,0.0,6.67,0.0,95.6,1,0,92270
2070,0,0,0,0,49,1,1,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),59.75,2934.3,1,40,33,35.87,6006,1,Seeley,0,0,DSL,32.790282,-115.689559,0,62.14,0,0,Offer B,1632,0,0,0,0,49,5,968.0,1757.63,0.0,2934.3,0,0,92273
2071,0,0,1,1,67,1,1,Fiber optic,0,1,1,0,Two year,0,Credit card (automatic),94.1,6302.8,0,53,27,11.4,4803,0,Thermal,0,0,Fiber Optic,33.53604,-116.119222,1,94.1,3,1,Offer A,17018,1,0,1,0,67,2,0.0,763.8000000000002,0.0,6302.8,0,1,92274
2072,1,0,0,1,39,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.35,779.2,0,42,0,48.61,2607,0,Salton City,0,1,NA,33.28156,-115.955541,0,19.35,0,0,None,799,0,0,0,0,39,1,0.0,1895.79,0.0,779.2,0,0,92275
2073,1,0,0,0,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,283.75,0,27,0,43.5,3854,0,Thousand Palms,0,1,NA,33.849263,-116.382778,0,19.9,0,0,Offer D,6242,0,0,0,0,14,1,0.0,609.0,0.0,283.75,1,0,92276
2074,0,1,0,0,43,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),108.15,4600.7,1,67,11,31.83,2833,1,Escondido,0,0,Cable,33.141265000000004,-116.967221,0,112.476,0,0,None,48690,1,0,0,0,43,2,506.0,1368.6899999999996,0.0,4600.7,0,0,92027
2075,1,1,0,0,56,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.05,5594,0,76,16,5.19,5514,0,Twentynine Palms,1,1,DSL,34.457829,-116.13958899999999,0,101.05,0,0,None,14104,0,0,0,0,56,1,0.0,290.6400000000001,0.0,5594.0,0,1,92278
2076,0,0,0,0,14,1,0,DSL,0,0,0,1,One year,0,Credit card (automatic),59.1,772.85,0,19,69,34.01,5718,0,Escondido,0,0,Cable,33.141265000000004,-116.967221,0,59.1,0,0,Offer D,48690,1,0,0,1,14,0,0.0,476.14,0.0,772.85,1,1,92027
2077,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,71.35,71.35,1,43,14,40.4,2619,1,Westmorland,0,0,DSL,33.03679,-115.60503,0,74.204,0,0,None,2388,0,1,0,0,1,6,0.0,40.4,0.0,71.35,0,1,92281
2078,1,0,1,1,16,1,0,DSL,1,1,0,0,One year,1,Mailed check,55.85,857.8,0,57,17,21.04,2464,0,White Water,0,1,DSL,33.972293,-116.654195,1,55.85,0,1,Offer D,805,0,0,1,0,16,2,146.0,336.64,0.0,857.8,0,0,92282
2079,1,0,1,1,70,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,106.05,7554.05,0,40,13,40.28,4583,0,Winterhaven,0,1,DSL,32.852947,-114.850784,1,106.05,1,1,Offer A,3663,0,0,1,1,70,0,0.0,2819.6,0.0,7554.05,0,1,92283
2080,1,1,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),84.1,5981.65,0,79,23,17.3,4671,0,Yucca Valley,1,1,Fiber Optic,34.159534,-116.42598400000001,1,84.1,0,1,None,20486,0,1,1,0,72,2,0.0,1245.6,0.0,5981.65,0,1,92284
2081,0,0,1,1,23,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.3,1702.9,0,51,75,48.73,5903,0,Landers,1,0,DSL,34.341737,-116.53941599999999,1,75.3,3,6,Offer D,2182,0,0,1,0,23,1,127.72,1120.79,0.0,1702.9,0,1,92285
2082,1,0,0,1,21,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,24.7,467.15,0,53,0,31.26,5403,0,Adelanto,0,1,NA,34.667815000000004,-117.53618300000001,0,24.7,1,0,Offer D,18980,0,0,0,0,21,0,0.0,656.46,0.0,467.15,0,0,92301
2083,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.15,20.15,1,42,0,21.59,4939,1,Amboy,0,0,NA,34.559882,-115.63716399999998,0,20.15,0,0,Offer E,42,0,0,0,0,1,4,0.0,21.59,0.0,20.15,0,0,92304
2084,1,0,0,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),69.75,69.75,1,35,20,27.97,2901,1,Angelus Oaks,0,1,Cable,34.1678,-116.86433000000001,0,72.54,0,0,Offer E,301,0,1,0,0,1,5,0.0,27.97,0.0,69.75,0,0,92305
2085,0,1,1,0,32,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.2,2931,1,69,7,33.74,5247,1,Fallbrook,0,0,DSL,33.362575,-117.299644,1,96.928,0,1,None,42239,0,0,1,0,32,5,205.0,1079.68,17.88,2931.0,0,0,92028
2086,1,0,1,1,17,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,80.85,1400.85,1,41,3,16.61,5174,1,Apple Valley,0,1,Fiber Optic,34.424926,-117.184503,1,84.084,0,1,None,28819,0,0,1,0,17,0,0.0,282.37,0.0,1400.85,0,1,92308
2087,0,0,0,0,4,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Electronic check,33.65,137.85,1,47,4,0.0,2563,1,Baker,0,0,Cable,35.28952,-116.09221399999998,0,34.996,0,0,Offer E,904,0,2,0,0,4,6,6.0,0.0,0.0,137.85,0,0,92309
2088,0,0,0,0,36,1,1,DSL,0,0,0,0,One year,0,Electronic check,55.8,1941.5,0,38,5,46.92,4770,0,Fort Irwin,1,0,DSL,35.349241,-116.77028100000001,0,55.8,0,0,None,9465,0,0,0,0,36,3,0.0,1689.12,0.0,1941.5,0,1,92310
2089,0,0,0,0,50,0,No phone service,DSL,0,1,0,0,Two year,0,Credit card (automatic),39.7,1932.75,0,48,6,0.0,5174,0,Barstow,1,0,DSL,34.965648,-117.00150900000001,0,39.7,0,0,None,31293,1,0,0,0,50,3,0.0,0.0,0.0,1932.75,0,1,92311
2090,0,0,1,1,48,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),29.5,1423.05,0,38,16,0.0,3194,0,Grand Terrace,0,0,Fiber Optic,34.029175,-117.30721100000001,1,29.5,1,6,None,11024,1,0,1,0,48,1,228.0,0.0,0.0,1423.05,0,0,92313
2091,0,0,0,1,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.15,970.85,0,40,0,18.95,4263,0,Big Bear City,0,0,NA,34.278967,-116.773825,0,20.15,3,0,None,9899,0,0,0,0,50,1,0.0,947.5,0.0,970.85,0,0,92314
2092,1,0,1,0,72,1,1,DSL,1,1,0,1,Two year,0,Credit card (automatic),79.55,5810.9,0,34,9,45.05,4766,0,Big Bear Lake,1,1,Cable,34.242058,-116.89801999999999,1,79.55,0,3,Offer A,5447,1,0,1,1,72,1,0.0,3243.6,0.0,5810.9,0,1,92315
2093,1,0,0,1,10,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),24.8,223.9,0,61,0,34.47,5212,0,Bloomington,0,1,NA,34.059722,-117.39103999999999,0,24.8,3,0,Offer D,25995,0,0,0,0,10,0,0.0,344.7,0.0,223.9,0,0,92316
2094,0,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,391.7,0,44,0,18.2,4333,0,Calimesa,0,0,NA,33.982787,-117.057627,0,19.65,0,0,Offer D,7334,0,0,0,0,18,2,0.0,327.6,0.0,391.7,0,0,92320
2095,1,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.95,79.95,1,56,6,3.13,4815,1,Cedar Glen,0,1,Cable,34.255203,-117.17565400000001,0,83.14800000000002,0,0,Offer E,455,0,0,0,0,1,3,0.0,3.13,0.0,79.95,0,0,92321
2096,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.3,19.3,1,58,0,25.62,3236,1,Colton,0,0,NA,34.030915,-117.273201,0,19.3,0,0,Offer E,52202,0,0,0,0,1,1,0.0,25.62,0.0,19.3,0,0,92324
2097,1,0,0,0,9,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.05,811.65,0,40,14,15.53,3475,0,Crestline,1,1,DSL,34.248061,-117.29028000000001,0,94.05,0,0,Offer E,10484,0,0,0,1,9,1,11.36,139.76999999999998,0.0,811.65,0,1,92325
2098,1,0,0,0,2,1,1,Fiber optic,1,0,0,1,Month-to-month,0,Mailed check,90.75,174.75,0,55,23,27.17,4766,0,Daggett,0,1,Fiber Optic,34.875144,-116.821698,0,90.75,0,0,Offer E,678,0,0,0,1,2,0,40.0,54.34,0.0,174.75,0,0,92327
2099,0,0,1,0,40,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),78.85,3126.85,0,61,17,39.97,5257,0,Death Valley,0,0,DSL,36.27688,-117.033326,1,78.85,0,10,None,443,1,0,1,0,40,0,532.0,1598.8,0.0,3126.85,0,0,92328
2100,1,0,1,0,69,1,1,Fiber optic,0,0,1,1,One year,0,Bank transfer (automatic),99.5,6841.45,0,50,4,3.81,4237,0,Essex,1,1,Cable,34.9436,-115.287901,1,99.5,0,10,Offer A,115,0,0,1,1,69,1,27.37,262.89,0.0,6841.45,0,1,92332
2101,0,0,1,0,37,1,1,Fiber optic,1,0,0,1,One year,1,Electronic check,99.2,3754.6,1,55,4,30.16,3599,1,Fawnskin,1,0,DSL,34.274846000000004,-116.93758100000001,1,103.16799999999999,0,1,None,414,1,2,1,1,37,4,150.0,1115.92,0.0,3754.6,0,0,92333
2102,1,0,0,1,18,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),80.55,1406.65,0,29,48,41.08,5334,0,Fontana,1,1,Fiber Optic,34.087558,-117.464096,0,80.55,3,0,Offer D,82630,0,0,0,0,18,1,0.0,739.4399999999998,0.0,1406.65,1,1,92335
2103,1,1,1,0,11,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.2,834.7,0,76,29,24.42,2848,0,Fontana,0,1,Fiber Optic,34.136367,-117.460803,1,70.2,0,7,Offer D,54586,0,0,1,0,11,0,24.21,268.62,0.0,834.7,0,1,92336
2104,0,0,1,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),85.2,627.4,1,32,18,26.41,2887,1,Fontana,0,0,DSL,34.049671000000004,-117.468896,1,88.60799999999999,0,0,Offer E,29847,0,2,0,1,8,1,113.0,211.28,0.0,627.4,0,0,92337
2105,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.25,242,1,40,28,17.87,5898,1,Ludlow,0,0,Fiber Optic,34.702766,-116.093376,0,78.26,0,0,None,23,0,0,0,0,3,3,68.0,53.61,0.0,242.0,0,0,92338
2106,1,0,1,1,55,1,0,DSL,1,0,0,1,One year,0,Credit card (automatic),59.45,3157,0,24,69,36.17,5712,0,Forest Falls,0,1,DSL,34.067699,-116.90389099999999,1,59.45,0,5,None,958,0,0,1,1,55,0,2178.0,1989.35,0.0,3157.0,1,0,92339
2107,1,0,1,0,33,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,93.35,3092,0,35,7,31.76,3348,0,Green Valley Lake,1,1,Cable,34.244411,-117.072654,1,93.35,0,5,None,317,0,1,1,1,33,1,0.0,1048.0800000000004,0.0,3092.0,0,1,92341
2108,0,0,0,0,46,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),44.95,2168.9,0,19,51,40.32,2626,0,Helendale,0,0,Cable,34.757783,-117.33997,0,44.95,0,0,None,4948,0,0,0,0,46,2,110.61,1854.72,0.0,2168.9,1,1,92342
2109,1,0,0,0,34,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),26.1,980.35,0,54,0,20.47,2026,0,Hesperia,0,1,NA,34.361387,-117.33750900000001,0,26.1,0,0,None,68515,0,0,0,0,34,0,0.0,695.98,0.0,980.35,0,0,92345
2110,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.2,65.95,0,64,0,31.81,4369,0,Highland,0,0,NA,34.129677,-117.15427700000001,0,20.2,0,0,None,48245,0,0,0,0,3,0,0.0,95.43,0.0,65.95,0,0,92346
2111,1,0,1,1,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,21.25,711.9,0,58,0,40.0,3047,0,Hinkley,0,1,NA,34.983808,-117.239306,1,21.25,3,6,None,1933,0,0,1,0,30,0,0.0,1200.0,0.0,711.9,0,0,92347
2112,0,0,0,0,33,1,1,DSL,1,0,0,0,One year,0,Electronic check,59.4,1952.8,0,41,7,10.28,2853,0,Lake Arrowhead,0,0,Cable,34.2565,-117.19335,0,59.4,0,0,None,9793,1,0,0,0,33,1,137.0,339.2399999999999,0.0,1952.8,0,0,92352
2113,1,0,1,1,45,1,1,Fiber optic,0,1,0,1,One year,1,Credit card (automatic),95.0,4368.85,0,25,69,33.45,2719,0,Loma Linda,1,1,Fiber Optic,34.049315,-117.255974,1,95.0,2,6,None,18068,0,0,1,1,45,0,3015.0,1505.2500000000002,0.0,4368.85,1,0,92354
2114,1,0,0,0,40,1,0,DSL,1,1,0,0,Month-to-month,1,Mailed check,61.9,2647.1,0,49,21,36.98,2520,0,Lucerne Valley,0,1,DSL,34.508417,-116.856103,0,61.9,0,0,None,5256,1,0,0,0,40,0,0.0,1479.1999999999996,0.0,2647.1,0,1,92356
2115,0,0,0,0,71,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,118.65,8477.6,0,58,21,17.9,4296,0,Lytle Creek,1,0,Fiber Optic,34.238162,-117.534306,0,118.65,0,0,Offer A,1090,1,0,0,1,71,2,1780.0,1270.9,0.0,8477.6,0,0,92358
2116,1,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,54.35,54.35,1,30,57,25.39,4212,1,Mentone,1,1,Cable,34.103578000000006,-117.04054,0,56.523999999999994,0,0,Offer E,7324,0,0,0,0,1,1,0.0,25.39,0.0,54.35,0,1,92359
2117,0,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),64.45,4528,0,53,6,0.0,5265,0,Needles,1,0,DSL,34.711224,-114.702256,1,64.45,0,0,Offer A,5488,1,0,0,1,72,2,27.17,0.0,0.0,4528.0,0,1,92363
2118,0,0,1,1,22,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.15,1790.65,0,59,29,33.46,4732,0,Nipton,0,0,Cable,35.478736,-115.51698400000001,1,80.15,3,5,Offer D,162,0,0,1,1,22,1,519.0,736.12,0.0,1790.65,0,0,92364
2119,1,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.2,845.6,0,44,0,4.72,2325,0,Temecula,0,1,NA,33.507255,-117.029473,1,20.2,0,6,None,46171,0,0,1,0,46,0,0.0,217.12,0.0,845.6,0,0,92592
2120,0,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,21.0,1210.3,0,53,0,38.51,5046,0,Oro Grande,0,0,NA,34.647959,-117.296957,1,21.0,3,8,Offer B,909,0,0,1,0,55,1,0.0,2118.05,0.0,1210.3,0,0,92368
2121,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.45,20.45,0,26,0,30.09,4845,0,Phelan,0,1,NA,34.441123,-117.53788600000001,0,20.45,0,0,None,12463,0,1,0,0,1,1,0.0,30.09,0.0,20.45,1,0,92371
2122,0,0,0,0,12,1,1,DSL,0,0,1,1,One year,1,Mailed check,75.85,854.45,0,23,47,49.25,5942,0,Pinon Hills,0,0,DSL,34.459322,-117.629729,0,75.85,0,0,Offer D,4280,1,0,0,1,12,0,0.0,591.0,0.0,854.45,1,1,92372
2123,1,0,0,0,31,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.45,2429.1,0,43,23,37.07,4684,0,Redlands,0,1,Fiber Optic,34.003243,-117.13828600000001,0,80.45,0,0,None,31230,0,0,0,0,31,0,0.0,1149.17,0.0,2429.1,0,1,92373
2124,1,0,1,0,5,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.95,100.4,1,37,8,0.0,5865,1,Redlands,0,1,Fiber Optic,34.064073,-117.16615800000001,1,25.948,0,1,Offer E,36675,0,1,1,0,5,3,8.0,0.0,0.0,100.4,0,0,92374
2125,0,0,1,1,67,1,1,DSL,1,0,1,1,Two year,1,Electronic check,75.5,5229.45,0,24,82,1.36,5420,0,Rialto,0,0,DSL,34.109775,-117.378904,1,75.5,0,5,Offer A,75882,0,0,1,1,67,0,4288.0,91.12,0.0,5229.45,1,0,92376
2126,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.45,44.45,0,45,16,23.34,3498,0,Rialto,0,1,DSL,34.156758,-117.40468600000001,0,44.45,0,0,None,18518,0,0,0,0,1,1,0.0,23.34,0.0,44.45,0,0,92377
2127,1,0,1,0,40,0,No phone service,DSL,1,1,0,0,One year,1,Electronic check,42.35,1716.45,1,39,23,0.0,5422,1,Running Springs,1,1,Cable,34.186211,-117.07683,1,44.044,0,1,Offer B,5395,0,0,1,0,40,7,395.0,0.0,0.0,1716.45,0,0,92382
2128,1,0,1,1,41,1,1,DSL,1,1,1,0,Month-to-month,1,Credit card (automatic),74.55,3023.55,0,61,20,28.55,2748,0,Shoshone,1,1,Fiber Optic,35.924252,-116.18866799999999,1,74.55,2,4,Offer B,87,0,0,1,0,41,1,0.0,1170.55,0.0,3023.55,0,1,92384
2129,1,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.3,75.3,1,38,20,39.44,3596,1,Sugarloaf,0,1,Cable,34.243088,-116.83001499999999,0,78.312,0,0,Offer E,1834,0,1,0,0,1,1,0.0,39.44,0.0,75.3,0,0,92386
2130,1,0,0,0,51,1,1,Fiber optic,1,1,1,0,One year,1,Electronic check,94.8,4837.6,1,22,64,44.77,5074,1,Fallbrook,0,1,Cable,33.362575,-117.299644,0,98.59200000000001,0,0,Offer B,42239,0,0,0,1,51,1,3096.0,2283.27,0.0,4837.6,1,0,92028
2131,1,0,1,1,42,0,No phone service,DSL,1,0,1,0,Two year,0,Credit card (automatic),48.15,2032.3,0,48,8,0.0,2673,0,Victorville,1,1,Fiber Optic,34.486835,-117.362274,1,48.15,0,10,Offer B,63235,1,0,1,0,42,1,163.0,0.0,0.0,2032.3,0,0,92392
2132,1,0,1,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.65,436.9,0,62,0,24.88,5460,0,Victorville,0,1,NA,34.567058,-117.362329,1,19.65,0,2,Offer D,12083,0,0,1,0,23,2,0.0,572.24,0.0,436.9,0,0,92394
2133,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.55,70.55,1,72,14,18.2,2146,1,Wrightwood,0,0,Cable,34.358321000000004,-117.61826299999998,0,73.372,0,0,Offer E,4253,0,0,0,0,1,4,0.0,18.2,0.0,70.55,0,0,92397
2134,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.15,20.15,0,40,0,27.59,3167,0,Yermo,0,0,NA,35.013298999999996,-116.834092,0,20.15,0,0,None,1195,0,0,0,0,1,0,0.0,27.59,0.0,20.15,0,0,92398
2135,0,0,0,0,56,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),106.6,5893.95,0,25,51,24.77,5056,0,Yucaipa,0,0,Fiber Optic,34.045970000000004,-117.011825,0,106.6,0,0,Offer B,41575,0,0,0,1,56,1,0.0,1387.12,0.0,5893.95,1,1,92399
2136,1,0,0,1,15,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,91.0,1430.05,0,31,12,30.22,4602,0,San Bernardino,0,1,Fiber Optic,34.105934999999995,-117.2914,0,91.0,1,0,Offer D,1779,0,0,0,0,15,3,17.16,453.3,0.0,1430.05,0,1,92401
2137,1,0,1,1,12,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.4,313,0,55,0,44.12,2219,0,San Bernardino,0,1,NA,34.183285999999995,-117.221722,1,25.4,3,8,Offer D,53636,0,0,1,0,12,0,0.0,529.4399999999998,0.0,313.0,0,0,92404
2138,0,0,1,1,54,1,0,DSL,1,0,0,1,Two year,0,Bank transfer (automatic),69.95,3871.85,0,21,76,28.17,5077,0,San Bernardino,1,0,Fiber Optic,34.142747,-117.30086399999999,1,69.95,0,3,Offer B,24644,1,0,1,1,54,1,2943.0,1521.18,0.0,3871.85,1,0,92405
2139,0,0,0,0,7,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,66.85,458.1,0,30,85,48.16,4858,0,San Bernardino,0,0,Fiber Optic,34.250069,-117.39394899999999,0,66.85,0,0,None,49355,0,1,0,1,7,1,0.0,337.12,0.0,458.1,0,1,92407
2140,0,0,1,1,33,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Credit card (automatic),86.15,2745.7,1,63,31,14.34,3336,1,San Bernardino,0,0,Cable,34.084909,-117.25810700000001,1,89.596,0,1,None,12149,0,1,1,1,33,3,851.0,473.22,0.0,2745.7,0,0,92408
2141,1,0,1,1,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.15,341.35,0,30,0,38.55,5271,0,San Bernardino,0,1,NA,34.106922,-117.29755300000001,1,20.15,3,4,Offer D,44556,0,1,1,0,16,1,0.0,616.8,0.0,341.35,0,0,92410
2142,0,0,0,1,21,1,0,DSL,1,0,0,1,One year,0,Mailed check,64.85,1336.8,0,55,15,30.88,3302,0,San Bernardino,1,0,DSL,34.122501,-117.32013799999999,0,64.85,0,0,Offer D,23146,0,0,0,1,21,2,0.0,648.48,0.0,1336.8,0,1,92411
2143,1,1,1,0,30,1,1,DSL,0,0,1,1,Two year,0,Electronic check,74.85,2181.75,0,77,8,40.5,5610,0,Riverside,1,1,DSL,33.994676,-117.372498,1,74.85,0,7,None,18999,0,0,1,0,30,0,175.0,1215.0,0.0,2181.75,0,0,92501
2144,1,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.5,147.75,0,45,25,26.38,5258,0,Riverside,0,1,DSL,33.890046000000005,-117.455583,0,50.5,0,0,None,71678,1,0,0,0,3,0,37.0,79.14,0.0,147.75,0,0,92503
2145,1,0,0,0,11,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,72.9,818.45,0,27,76,18.33,3042,0,Riverside,1,1,Cable,33.9108,-117.39815300000001,0,72.9,0,0,Offer D,46550,0,0,0,0,11,0,0.0,201.63,0.0,818.45,1,1,92504
2146,0,0,0,0,62,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),115.05,7133.45,0,39,13,36.84,6494,0,Riverside,1,0,DSL,33.920907,-117.489426,0,115.05,0,0,Offer B,38446,1,0,0,1,62,0,0.0,2284.080000000001,0.0,7133.45,0,1,92505
2147,1,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.0,348.8,0,42,0,33.16,5379,0,Riverside,0,1,NA,33.930931,-117.36178799999999,0,19.0,0,0,Offer D,42425,0,2,0,0,18,1,0.0,596.8799999999999,0.0,348.8,0,0,92506
2148,1,0,0,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.55,128.6,0,20,0,17.53,2309,0,Riverside,0,1,NA,33.976328,-117.31978600000001,0,19.55,1,0,None,48649,0,1,0,0,6,1,0.0,105.18,0.0,128.6,1,0,92507
2149,0,0,0,0,46,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,101.1,4674.4,0,45,22,27.97,4883,0,Riverside,1,0,DSL,33.885498999999996,-117.324959,0,101.1,0,0,Offer B,17147,0,0,0,1,46,3,0.0,1286.62,0.0,4674.4,0,1,92508
2150,1,0,0,0,21,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.1,1737.45,0,46,9,49.05,4649,0,Riverside,0,1,Cable,34.004379,-117.447864,0,84.1,0,0,None,63999,0,0,0,1,21,0,15.64,1030.05,0.0,1737.45,0,1,92509
2151,1,0,0,0,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.15,1498.85,0,45,0,37.79,5987,0,March Air Reserve Base,0,1,NA,33.888323,-117.277533,0,24.15,0,0,None,1005,0,0,0,0,68,0,0.0,2569.72,0.0,1498.85,0,0,92518
2152,0,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.1,50.1,0,19,51,29.13,5617,0,Lake Elsinore,0,0,DSL,33.655421000000004,-117.391751,0,50.1,0,0,None,38519,0,0,0,0,1,2,0.0,29.13,0.0,50.1,1,0,92530
2153,0,0,1,0,25,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.6,1797.75,0,26,82,37.1,4591,0,Lake Elsinore,1,0,Fiber Optic,33.705836,-117.31820400000001,1,74.6,0,7,None,4546,0,0,1,0,25,0,0.0,927.5,0.0,1797.75,1,1,92532
2154,0,0,0,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,498.1,0,57,0,34.24,2639,0,Aguanga,0,0,NA,33.482243,-116.827173,0,19.75,1,0,None,2433,0,0,0,0,24,0,0.0,821.76,0.0,498.1,0,0,92536
2155,0,0,1,0,30,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.0,2624.25,1,25,45,4.82,3698,1,Anza,0,0,Cable,33.527605,-116.666551,1,88.4,0,1,Offer C,3745,0,0,1,1,30,2,1181.0,144.60000000000005,0.0,2624.25,1,0,92539
2156,0,0,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,80.55,184.1,1,29,45,33.89,2856,1,Hemet,0,0,Fiber Optic,33.739415,-116.96833899999999,0,83.772,0,0,Offer E,29687,0,0,0,1,2,5,83.0,67.78,0.0,184.1,1,0,92543
2157,1,0,1,0,51,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),106.8,5498.8,0,31,21,29.4,4640,0,Hemet,1,1,Fiber Optic,33.644585,-116.871544,1,106.8,0,3,Offer B,39264,0,0,1,1,51,0,115.47,1499.4,0.0,5498.8,0,1,92544
2158,0,0,1,1,57,1,1,DSL,1,0,1,1,Two year,1,Electronic check,84.5,4845.4,0,33,16,10.05,5928,0,Hemet,1,0,Fiber Optic,33.734933000000005,-117.044145,1,84.5,0,2,Offer B,25694,1,0,1,1,57,1,0.0,572.85,0.0,4845.4,0,1,92545
2159,0,0,0,0,15,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.05,369.1,0,52,0,40.97,5218,0,Homeland,0,0,NA,33.761894,-117.12086799999999,0,25.05,0,0,None,4283,0,2,0,0,15,2,0.0,614.55,0.0,369.1,0,0,92548
2160,0,0,1,1,72,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),83.7,6096.9,0,25,46,16.05,4592,0,Idyllwild,1,0,DSL,33.755039000000004,-116.741796,1,83.7,0,9,None,3588,1,0,1,1,72,0,0.0,1155.6,0.0,6096.9,1,1,92549
2161,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.8,160.75,1,37,18,24.31,5270,1,Moreno Valley,1,0,Cable,33.882740000000005,-117.224878,0,78.832,0,0,Offer E,22983,0,0,0,0,2,0,29.0,48.62,0.0,160.75,0,0,92551
2162,1,0,1,0,28,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Credit card (automatic),96.6,2684.35,0,25,52,33.57,5530,0,Moreno Valley,1,1,Fiber Optic,33.923149,-117.244933,1,96.6,0,10,None,61205,0,0,1,0,28,0,139.59,939.96,0.0,2684.35,1,1,92553
2163,1,1,1,0,29,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.5,3004.15,1,75,31,25.78,5137,1,Moreno Valley,1,1,Fiber Optic,33.907361,-117.109972,1,102.44,0,1,None,12743,0,0,1,1,29,4,931.0,747.62,37.55,3004.15,0,0,92555
2164,1,0,1,1,70,1,0,Fiber optic,1,1,1,0,Two year,1,Credit card (automatic),101.1,6994.8,0,52,19,49.67,4226,0,Moreno Valley,1,1,Fiber Optic,33.970661,-117.255039,1,101.1,2,10,None,46214,1,0,1,0,70,0,132.9,3476.9,0.0,6994.8,0,1,92557
2165,0,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.2,273.25,0,52,0,26.57,2953,0,Mountain Center,0,0,NA,33.638645000000004,-116.55783000000001,0,20.2,0,0,None,1500,0,0,0,0,13,1,0.0,345.41,0.0,273.25,0,0,92561
2166,0,1,1,0,59,1,1,Fiber optic,1,1,0,0,One year,1,Electronic check,94.05,5483.9,0,71,13,19.14,5061,0,Murrieta,1,0,Cable,33.548869,-117.33416499999998,1,94.05,0,0,None,36149,1,0,0,0,59,0,713.0,1129.26,0.0,5483.9,0,0,92562
2167,1,1,1,0,13,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.25,1233.65,1,67,7,31.7,2982,1,Murrieta,0,1,Fiber Optic,33.581045,-117.14719,1,99.06,0,1,None,18311,0,2,1,1,13,3,86.0,412.1,48.09,1233.65,0,0,92563
2168,1,1,1,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.4,527.9,1,72,19,8.92,4969,1,Nuevo,0,1,DSL,33.827690000000004,-117.102244,1,77.376,0,1,None,7344,0,0,1,0,7,5,0.0,62.44,32.46,527.9,0,1,92567
2169,0,0,1,0,62,1,0,DSL,1,0,1,1,Two year,0,Mailed check,81.0,4985.9,0,49,22,13.32,4684,0,Perris,1,0,DSL,33.787298,-117.320676,1,81.0,0,6,Offer B,36817,1,0,1,1,62,0,1097.0,825.84,0.0,4985.9,0,0,92570
2170,0,0,0,0,21,1,0,DSL,1,0,0,0,One year,1,Electronic check,60.25,1258.35,0,30,51,7.41,4870,0,Perris,1,0,DSL,33.828289,-117.20166599999999,0,60.25,0,0,None,26357,1,0,0,0,21,0,64.18,155.61,0.0,1258.35,0,1,92571
2171,0,0,0,0,2,1,0,DSL,0,0,0,1,Month-to-month,0,Electronic check,60.85,111.4,0,28,82,15.25,3796,0,San Jacinto,1,0,DSL,33.806708,-117.02006999999999,0,60.85,0,0,None,4456,0,0,0,1,2,1,91.0,30.5,0.0,111.4,1,0,92582
2172,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),43.95,43.95,0,38,5,45.59,5684,0,San Jacinto,0,0,DSL,33.796568,-116.924723,0,43.95,0,0,None,21349,0,0,0,0,1,2,0.0,45.59,0.0,43.95,0,1,92583
2173,1,0,0,0,4,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,86.05,308.1,0,63,20,44.36,3653,0,Menifee,1,1,Cable,33.653338,-117.178271,0,86.05,0,0,None,14068,0,0,0,1,4,2,0.0,177.44,0.0,308.1,0,1,92584
2174,0,0,0,0,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.25,383.65,0,45,0,18.57,5586,0,Sun City,0,0,NA,33.739412,-117.17333400000001,0,20.25,0,0,None,8692,0,0,0,0,19,0,0.0,352.83,0.0,383.65,0,0,92585
2175,0,0,0,0,30,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,85.15,2555.9,1,45,9,9.34,4417,1,Sun City,0,0,Cable,33.707483,-117.200006,0,88.55600000000003,0,0,Offer C,18161,1,1,0,0,30,4,230.0,280.2,0.0,2555.9,0,0,92586
2176,1,0,1,1,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.4,1284.2,0,48,0,5.48,4890,0,Sun City,0,1,NA,33.69887,-117.25071000000001,1,19.4,2,6,None,13151,0,0,1,0,67,0,0.0,367.16,0.0,1284.2,0,0,92587
2177,1,1,1,0,72,1,1,Fiber optic,1,1,0,1,Two year,1,Credit card (automatic),102.65,7550.3,0,75,5,28.5,4680,0,Temecula,1,1,Fiber Optic,33.475493,-117.219551,1,102.65,0,5,None,3070,0,0,1,0,72,1,378.0,2052.0,0.0,7550.3,0,0,92590
2178,1,0,1,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.9,1110.05,0,35,0,34.46,4157,0,Temecula,0,1,NA,33.540603999999995,-117.10909,1,19.9,0,8,Offer B,25655,0,0,1,0,53,0,0.0,1826.38,0.0,1110.05,0,0,92591
2179,0,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.55,99.6,0,54,0,37.97,2575,0,Temecula,0,0,NA,33.507255,-117.029473,0,19.55,0,0,None,46171,0,0,0,0,5,1,0.0,189.85,0.0,99.6,0,0,92592
2180,1,1,1,0,71,1,0,Fiber optic,0,1,0,1,Two year,1,Credit card (automatic),95.5,6707.15,0,75,9,1.23,6412,0,Wildomar,1,1,Cable,33.617108,-117.253349,1,95.5,0,2,None,19368,1,0,1,0,71,0,0.0,87.33,0.0,6707.15,0,1,92595
2181,0,0,1,1,50,1,1,DSL,0,1,1,1,One year,1,Credit card (automatic),84.15,4164.4,0,53,11,46.49,4625,0,Winchester,1,0,Fiber Optic,33.657433000000005,-117.04253999999999,1,84.15,0,9,Offer B,4093,1,0,1,1,50,2,458.0,2324.5,0.0,4164.4,0,0,92596
2182,1,0,1,1,56,1,1,Fiber optic,0,0,1,1,Two year,1,Electronic check,103.2,5873.75,0,38,19,42.16,4478,0,Irvine,1,1,DSL,33.720359,-117.733655,1,103.2,1,3,Offer B,2762,1,0,1,1,56,2,0.0,2360.96,0.0,5873.75,0,1,92602
2183,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),50.2,109.25,0,61,28,6.34,4697,0,Irvine,0,1,Fiber Optic,33.688546,-117.788091,0,50.2,0,0,None,27369,1,0,0,0,2,1,31.0,12.68,0.0,109.25,0,0,92604
2184,0,1,0,0,2,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,88.55,179.25,1,68,31,21.57,3685,1,Irvine,1,0,Cable,33.703976000000004,-117.82417199999999,0,92.09200000000001,0,0,None,17621,0,6,0,1,2,3,56.0,43.14,0.0,179.25,0,0,92606
2185,1,0,1,1,24,1,1,DSL,1,0,0,0,Month-to-month,0,Electronic check,54.75,1338.15,1,63,20,17.27,5699,1,Foothill Ranch,0,1,Cable,33.698728,-117.67768000000001,1,56.94000000000001,2,1,Offer C,10936,0,0,1,0,24,6,268.0,414.48,0.0,1338.15,0,0,92610
2186,1,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.95,862.4,0,40,0,26.12,3574,0,Irvine,0,1,NA,33.643095,-117.810896,1,19.95,2,9,Offer B,41062,0,0,1,0,46,2,0.0,1201.52,0.0,862.4,0,0,92612
2187,1,0,1,0,71,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,116.25,8564.75,0,42,9,6.19,6124,0,Irvine,1,1,Fiber Optic,33.680302000000005,-117.83329599999999,1,116.25,0,4,None,22499,1,0,1,1,71,0,0.0,439.49,0.0,8564.75,0,1,92614
2188,0,0,0,0,29,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,31.2,926.2,0,30,59,0.0,4761,0,Irvine,0,0,Fiber Optic,33.667145,-117.73213500000001,0,31.2,0,0,None,6301,1,0,0,0,29,0,54.65,0.0,0.0,926.2,0,1,92618
2189,1,0,1,1,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.45,1718.2,0,23,0,33.09,5295,0,Irvine,0,1,NA,33.716136,-117.752574,1,24.45,3,1,None,26419,0,0,1,0,69,1,0.0,2283.21,0.0,1718.2,1,0,92620
2190,1,0,1,0,71,1,1,DSL,0,1,1,1,Two year,0,Credit card (automatic),84.2,5956.85,0,32,30,15.12,4753,0,Capistrano Beach,1,1,Fiber Optic,33.458754,-117.665104,1,84.2,0,4,None,7465,1,0,1,1,71,2,0.0,1073.52,0.0,5956.85,0,1,92624
2191,0,1,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,91.3,91.3,1,68,2,43.61,2371,1,Corona Del Mar,0,0,Fiber Optic,33.600986999999996,-117.862734,0,94.95200000000001,0,0,None,13422,0,0,0,1,1,0,0.0,43.61,0.0,91.3,0,0,92625
2192,1,1,1,0,56,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),85.65,4824.45,0,71,30,31.68,6500,0,Costa Mesa,1,1,DSL,33.678591,-117.90547099999999,1,85.65,0,8,None,48207,1,0,1,0,56,0,1447.0,1774.08,0.0,4824.45,0,0,92626
2193,1,0,0,1,56,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,21.2,1238.65,0,38,0,48.63,6473,0,Costa Mesa,0,1,NA,33.645672,-117.92261299999998,0,21.2,0,0,Offer B,62069,0,0,0,0,56,1,0.0,2723.28,0.0,1238.65,0,0,92627
2194,1,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.5,79.5,1,60,25,48.97,4490,1,Dana Point,0,1,Cable,33.477923,-117.70531399999999,0,82.68,0,0,Offer E,27730,0,0,0,0,1,1,0.0,48.97,0.0,79.5,0,0,92629
2195,0,0,1,0,28,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,25.55,672.2,0,22,0,43.36,3493,0,Lake Forest,0,0,NA,33.644849,-117.68425400000001,1,25.55,0,7,None,59176,0,0,1,0,28,0,0.0,1214.08,0.0,672.2,1,0,92630
2196,0,0,1,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.2,382.2,0,47,0,46.91,3636,0,Huntington Beach,0,0,NA,33.666301000000004,-117.969501,1,20.2,2,6,None,56517,0,0,1,0,19,0,0.0,891.29,0.0,382.2,0,0,92646
2197,1,0,1,0,66,1,1,DSL,0,0,0,1,Month-to-month,0,Electronic check,63.85,4264.6,0,21,69,7.67,5956,0,Huntington Beach,0,1,Fiber Optic,33.723579,-118.00544099999999,1,63.85,0,4,None,58764,1,0,1,1,66,0,2943.0,506.22,0.0,4264.6,1,0,92647
2198,0,0,1,1,17,1,1,DSL,0,0,0,0,One year,1,Mailed check,61.95,1070.7,0,52,25,47.59,4759,0,Huntington Beach,1,0,DSL,33.679659,-118.016195,1,61.95,0,6,None,42663,1,2,1,0,17,3,26.77,809.0300000000002,0.0,1070.7,0,1,92648
2199,1,0,1,1,52,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.75,1345.85,0,61,0,49.51,4676,0,Huntington Beach,0,1,NA,33.721917,-118.043237,1,25.75,2,6,Offer B,32304,0,0,1,0,52,1,0.0,2574.52,0.0,1345.85,0,0,92649
2200,0,0,0,0,19,1,0,DSL,0,1,1,0,One year,0,Electronic check,58.2,1045.25,0,19,69,24.35,4033,0,Laguna Beach,0,0,Fiber Optic,33.570023,-117.773669,0,58.2,0,0,None,25206,0,0,0,0,19,1,721.0,462.65,0.0,1045.25,1,0,92651
2201,0,0,0,0,36,1,0,DSL,1,1,1,1,One year,0,Bank transfer (automatic),85.85,3003.55,0,26,73,13.9,4898,0,Laguna Hills,1,0,DSL,33.606899,-117.717854,0,85.85,0,0,None,48273,1,0,0,1,36,1,0.0,500.4,0.0,3003.55,1,1,92653
2202,1,1,1,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.1,467.55,1,75,24,16.05,3669,1,Midway City,0,1,DSL,33.744439,-117.98588000000001,1,72.904,0,1,None,8660,0,0,1,0,7,2,0.0,112.35,20.23,467.55,0,1,92655
2203,1,0,1,1,72,1,1,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),104.9,7537.5,0,22,52,41.18,4927,0,Aliso Viejo,1,1,Fiber Optic,33.571259000000005,-117.731917,1,104.9,2,9,None,41237,1,0,1,1,72,1,0.0,2964.96,0.0,7537.5,1,1,92656
2204,1,0,1,1,67,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,111.3,7482.1,1,58,23,29.24,4146,1,Newport Coast,1,1,Cable,33.603282,-117.82184099999999,1,115.75200000000001,0,0,Offer A,5597,0,0,0,1,67,3,1721.0,1959.08,0.0,7482.1,0,0,92657
2205,1,1,0,0,34,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,99.85,3343.15,0,72,12,35.0,5626,0,Newport Beach,1,1,DSL,33.634626000000004,-117.874882,0,99.85,0,0,None,28687,0,0,0,0,34,0,401.0,1190.0,0.0,3343.15,0,0,92660
2206,1,1,1,0,57,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),95.25,5427.05,1,74,23,49.91,6259,1,Newport Beach,1,1,Cable,33.601309,-117.902304,1,99.06,0,1,None,4242,0,0,1,0,57,5,1248.0,2844.87,12.59,5427.05,0,0,92661
2207,0,0,1,0,7,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.25,587.1,1,63,29,44.66,3344,1,Newport Beach,1,0,Cable,33.606336,-117.893042,1,89.7,0,1,Offer E,3124,0,0,1,0,7,1,170.0,312.62,0.0,587.1,0,0,92662
2208,0,1,1,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.8,100.8,1,78,25,17.35,3128,1,Newport Beach,1,0,Cable,33.62251,-117.927024,1,104.83200000000001,0,4,None,22133,0,1,1,0,1,2,0.0,17.35,0.0,100.8,0,0,92663
2209,1,0,1,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.55,161.15,0,38,0,22.34,4909,0,San Clemente,0,1,NA,33.429488,-117.60943200000001,1,19.55,0,7,None,34946,0,0,1,0,8,0,0.0,178.72,0.0,161.15,0,0,92672
2210,0,0,0,0,69,1,1,Fiber optic,0,0,1,1,Two year,0,Electronic check,104.0,7028.5,0,44,13,1.85,5902,0,San Clemente,1,0,DSL,33.4725,-117.584273,0,104.0,0,0,None,15297,1,0,0,1,69,0,914.0,127.65,0.0,7028.5,0,0,92673
2211,0,0,1,0,50,1,1,Fiber optic,1,0,1,1,One year,1,Mailed check,104.4,5232.9,0,57,7,20.79,6100,0,San Juan Capistrano,1,0,DSL,33.521446999999995,-117.60255500000001,1,104.4,0,7,Offer B,34321,0,0,1,1,50,0,366.0,1039.5,0.0,5232.9,0,0,92675
2212,1,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.5,225.85,0,58,0,15.71,5039,0,Silverado,0,1,NA,33.782346000000004,-117.635263,0,19.5,0,0,None,1859,0,0,0,0,10,1,0.0,157.10000000000005,0.0,225.85,0,0,92676
2213,0,0,1,1,12,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.25,274.7,0,39,0,39.59,2646,0,Laguna Niguel,0,0,NA,33.529047,-117.701175,1,25.25,2,4,None,62103,0,0,1,0,12,0,0.0,475.08,0.0,274.7,0,0,92677
2214,0,0,0,0,14,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,86.3,1180.95,1,64,29,29.3,3677,1,Trabuco Canyon,0,0,Fiber Optic,33.631119,-117.567346,0,89.75200000000001,0,0,None,32268,0,0,0,1,14,0,342.0,410.2,0.0,1180.95,0,0,92679
2215,0,0,1,0,70,0,No phone service,DSL,1,0,0,1,Two year,1,Bank transfer (automatic),49.85,3370.2,0,46,26,0.0,5460,0,Westminster,1,0,Fiber Optic,33.752590999999995,-117.99366100000002,1,49.85,0,8,None,88230,1,0,1,1,70,1,87.63,0.0,0.0,3370.2,0,1,92683
2216,0,1,0,0,64,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),108.95,7111.3,0,76,24,22.86,5780,0,Rancho Santa Margarita,1,0,DSL,33.624654,-117.611733,0,108.95,0,0,None,42193,1,0,0,0,64,1,1707.0,1463.04,0.0,7111.3,0,0,92688
2217,0,0,1,1,66,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.9,5958.85,0,31,3,36.36,4082,0,Mission Viejo,1,0,DSL,33.611945,-117.66586699999999,1,89.9,0,9,None,46371,1,0,1,1,66,2,17.88,2399.76,0.0,5958.85,0,1,92691
2218,0,0,1,1,71,1,0,DSL,1,0,1,1,Two year,1,Credit card (automatic),82.0,5999.85,0,40,23,38.22,5770,0,Mission Viejo,1,0,Fiber Optic,33.60693,-117.644253,1,82.0,0,0,None,46227,1,1,0,1,71,1,1380.0,2713.62,0.0,5999.85,0,0,92692
2219,1,1,0,0,20,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,89.95,1648.45,0,70,23,48.46,4812,0,Ladera Ranch,0,1,Fiber Optic,33.569186,-117.640055,0,89.95,0,0,Offer D,350,0,0,0,0,20,0,379.0,969.2,0.0,1648.45,0,0,92694
2220,1,0,1,0,72,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),79.35,5753.25,0,48,14,29.8,4278,0,Santa Ana,0,1,Fiber Optic,33.748478000000006,-117.85891799999999,1,79.35,0,2,None,58157,1,0,1,1,72,0,805.0,2145.6,0.0,5753.25,0,0,92701
2221,0,0,1,1,71,1,0,DSL,1,1,0,0,Two year,0,Credit card (automatic),64.05,4492.9,0,64,29,4.71,4374,0,Santa Ana,1,0,Fiber Optic,33.748635,-117.906125,1,64.05,0,10,None,70011,1,0,1,0,71,0,1303.0,334.41,0.0,4492.9,0,0,92703
2222,1,0,1,1,38,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),101.15,3956.7,0,34,14,24.22,3738,0,Santa Ana,1,1,Fiber Optic,33.719869,-117.907063,1,101.15,1,9,None,91188,0,0,1,1,38,0,554.0,920.36,0.0,3956.7,0,0,92704
2223,0,0,0,0,28,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.95,2625.55,1,56,33,30.28,2468,1,Santa Ana,0,0,DSL,33.766003999999995,-117.786763,0,93.54799999999999,0,0,Offer C,44117,0,1,0,1,28,6,866.0,847.84,0.0,2625.55,0,0,92705
2224,1,1,1,0,17,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,76.45,1233.4,1,66,9,1.05,3266,1,Santa Ana,0,1,Fiber Optic,33.765893,-117.881533,1,79.50800000000002,0,2,None,37879,0,3,1,0,17,5,111.0,17.85,0.0,1233.4,0,0,92706
2225,1,0,0,0,33,0,No phone service,DSL,0,1,1,0,One year,1,Electronic check,39.1,1309,0,62,30,0.0,2855,0,Santa Ana,0,1,Fiber Optic,33.714828999999995,-117.872941,0,39.1,0,0,None,62634,0,0,0,0,33,1,0.0,0.0,0.0,1309.0,0,1,92707
2226,0,0,1,1,23,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,34.6,813.45,0,27,42,0.0,4445,0,Fountain Valley,0,0,Fiber Optic,33.712036,-117.95011299999999,1,34.6,0,10,None,54548,1,0,1,0,23,0,342.0,0.0,0.0,813.45,1,0,92708
2227,1,0,1,1,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,19.55,1108.8,0,54,0,27.93,4801,0,Tustin,0,1,NA,33.735802,-117.818805,1,19.55,0,3,Offer B,55062,0,0,1,0,58,0,0.0,1619.94,0.0,1108.8,0,0,92780
2228,0,1,1,0,70,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),104.45,7349.35,0,73,13,39.34,5004,0,Tustin,0,0,DSL,33.738543,-117.785046,1,104.45,0,3,Offer A,17494,1,0,1,0,70,2,955.0,2753.8,0.0,7349.35,0,0,92782
2229,1,0,1,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.5,294.2,0,40,5,28.47,2896,0,Anaheim,0,1,DSL,33.844983,-117.952151,1,70.5,0,2,None,60553,0,0,1,0,4,0,0.0,113.88,0.0,294.2,0,1,92801
2230,1,0,1,1,45,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.35,929.2,0,24,0,39.03,4210,0,Anaheim,0,1,NA,33.807864,-117.923782,1,20.35,2,3,Offer B,45086,0,0,1,0,45,1,0.0,1756.35,0.0,929.2,1,0,92802
2231,1,0,0,0,10,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.0,740,1,41,30,27.28,3156,1,Anaheim,0,1,Cable,33.818000000000005,-117.974404,0,72.8,0,0,None,81333,0,1,0,0,10,2,222.0,272.8,0.0,740.0,0,0,92804
2232,1,0,1,1,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.45,754.5,0,26,0,32.3,5745,0,Anaheim,0,1,NA,33.830209,-117.906099,1,19.45,2,2,None,68802,0,0,1,0,36,1,0.0,1162.8,0.0,754.5,1,0,92805
2233,1,0,0,0,54,1,0,DSL,1,1,1,0,Month-to-month,1,Mailed check,69.9,3883.3,0,61,24,27.62,6092,0,Anaheim,0,1,DSL,33.837959999999995,-117.870494,0,69.9,0,0,Offer B,34398,1,0,0,0,54,0,0.0,1491.48,0.0,3883.3,0,1,92806
2234,1,0,1,1,23,1,1,DSL,0,1,0,0,Two year,0,Mailed check,59.7,1414.2,0,33,17,13.79,3464,0,Anaheim,0,1,Cable,33.848733,-117.788357,1,59.7,0,6,None,36301,1,0,1,0,23,0,240.0,317.17,0.0,1414.2,0,0,92807
2235,0,0,1,1,41,1,1,DSL,1,1,1,0,One year,1,Credit card (automatic),78.35,3211.2,0,28,26,18.84,2894,0,Anaheim,1,0,Fiber Optic,33.850452000000004,-117.72666799999999,1,78.35,0,8,Offer B,19629,0,0,1,0,41,1,0.0,772.4399999999998,0.0,3211.2,1,1,92808
2236,1,1,0,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,71.45,371.6,0,78,9,17.13,5171,0,Brea,0,1,Fiber Optic,33.930199,-117.862898,0,71.45,0,0,Offer E,34055,0,0,0,0,5,0,0.0,85.64999999999998,0.0,371.6,0,1,92821
2237,1,0,1,1,27,0,No phone service,DSL,0,1,0,1,One year,1,Credit card (automatic),45.85,1246.4,0,25,27,0.0,2068,0,Brea,1,1,Fiber Optic,33.924143,-117.79387,1,45.85,0,3,None,1408,0,0,1,1,27,1,337.0,0.0,0.0,1246.4,1,0,92823
2238,0,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.85,95.85,0,50,14,2.7,3270,0,Fullerton,0,0,Cable,33.879983,-117.895482,0,95.85,0,0,None,34592,1,0,0,1,1,0,0.0,2.7,0.0,95.85,0,1,92831
2239,0,0,1,1,67,0,No phone service,DSL,1,0,0,0,Two year,0,Credit card (automatic),35.7,2545.7,0,55,30,0.0,5655,0,Fullerton,0,0,Fiber Optic,33.868316,-117.929029,1,35.7,0,5,None,24502,1,0,1,0,67,0,0.0,0.0,0.0,2545.7,0,1,92832
2240,0,1,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),89.55,6448.85,0,74,24,5.77,4993,0,Fullerton,1,0,DSL,33.877639,-117.96121200000002,1,89.55,0,4,Offer A,46105,1,0,1,0,72,0,0.0,415.44,0.0,6448.85,0,1,92833
2241,0,0,1,1,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.95,1468.9,0,40,0,29.06,5243,0,Fullerton,0,0,NA,33.902211,-117.914922,1,24.95,2,9,None,21157,0,0,1,0,56,2,0.0,1627.36,0.0,1468.9,0,0,92835
2242,1,0,1,1,44,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,24.85,1013.6,0,44,0,32.22,5331,0,Garden Grove,0,1,NA,33.787165,-117.93188899999998,1,24.85,0,7,None,50641,0,0,1,0,44,1,0.0,1417.6799999999996,0.0,1013.6,0,0,92840
2243,0,1,1,0,66,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.8,6690.75,0,73,20,28.06,5469,0,Garden Grove,0,0,DSL,33.786738,-117.982564,1,100.8,0,0,Offer A,31428,0,0,0,0,66,2,0.0,1851.96,0.0,6690.75,0,1,92841
2244,0,0,0,0,34,1,1,DSL,1,1,0,0,One year,1,Mailed check,64.4,2088.75,1,53,4,34.41,5189,1,Garden Grove,0,0,DSL,33.764018,-117.93150700000001,0,66.97600000000001,0,0,Offer C,43491,1,1,0,0,34,6,84.0,1169.9399999999996,0.0,2088.75,0,0,92843
2245,0,0,1,0,69,1,1,Fiber optic,0,0,1,1,Two year,0,Bank transfer (automatic),105.35,7240.65,0,51,6,14.69,5268,0,Garden Grove,1,0,Cable,33.766476000000004,-117.96979499999999,1,105.35,0,3,None,23481,1,2,1,1,69,1,434.0,1013.61,0.0,7240.65,0,0,92844
2246,0,0,1,1,1,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,102.45,102.45,1,52,10,25.88,4811,1,Garden Grove,1,0,Fiber Optic,33.782955,-118.02645600000001,1,106.54799999999999,0,1,None,15878,0,0,1,1,1,2,0.0,25.88,0.0,102.45,0,0,92845
2247,0,0,0,0,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.65,830.25,0,48,0,26.03,3878,0,Norco,0,0,NA,33.925833000000004,-117.55963899999999,0,19.65,0,0,None,22443,0,2,0,0,40,2,0.0,1041.2,0.0,830.25,0,0,92860
2248,1,0,1,1,30,1,1,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),54.45,1588.7,0,50,19,12.49,2613,0,Villa Park,0,1,Cable,33.817473,-117.81046200000002,1,54.45,2,6,None,5935,0,1,1,0,30,2,0.0,374.7,0.0,1588.7,0,1,92861
2249,0,0,0,0,11,1,0,DSL,0,0,1,1,Month-to-month,0,Mailed check,70.5,829.3,0,38,12,47.61,5541,0,Orange,0,0,DSL,33.828779,-117.848299,0,70.5,0,0,None,18058,1,0,0,1,11,0,9.95,523.71,0.0,829.3,0,1,92865
2250,0,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.1,302.45,0,58,0,9.74,4359,0,Orange,0,0,NA,33.784597,-117.84453500000001,0,20.1,0,0,None,15396,0,1,0,0,15,1,0.0,146.1,0.0,302.45,0,0,92866
2251,1,0,0,0,11,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,69.35,712.25,0,35,8,16.14,2288,0,Orange,1,1,Fiber Optic,33.81859,-117.821288,0,69.35,0,0,None,40915,0,0,0,1,11,0,57.0,177.54000000000005,0.0,712.25,0,0,92867
2252,0,0,1,1,64,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.8,1336.65,0,47,0,23.25,5384,0,Orange,0,0,NA,33.787796,-117.875928,1,19.8,0,7,None,23172,0,0,1,0,64,0,0.0,1488.0,0.0,1336.65,0,0,92868
2253,1,1,1,0,72,1,0,DSL,1,1,1,0,Two year,0,Bank transfer (automatic),74.4,5360.75,0,69,9,5.27,5590,0,Orange,1,1,Fiber Optic,33.792790999999994,-117.789749,1,74.4,0,7,Offer A,37916,1,0,1,0,72,3,482.0,379.44,0.0,5360.75,0,0,92869
2254,1,1,1,0,72,1,1,Fiber optic,1,1,0,0,Two year,1,Bank transfer (automatic),93.05,6735.05,0,73,30,1.34,4988,0,Placentia,1,1,DSL,33.881158,-117.85478300000001,1,93.05,0,10,Offer A,48170,1,0,1,0,72,0,2021.0,96.48,0.0,6735.05,0,0,92870
2255,0,0,0,1,1,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,51.2,51.2,0,42,26,2.98,3699,0,Corona,0,0,Fiber Optic,33.893823,-117.531446,0,51.2,3,0,None,44875,0,0,0,0,1,0,0.0,2.98,0.0,51.2,0,0,92879
2256,0,0,0,1,15,1,0,DSL,1,1,0,0,One year,0,Credit card (automatic),65.6,1010,0,26,73,20.11,2976,0,Corona,1,0,Fiber Optic,33.918043,-117.61780900000001,0,65.6,0,0,Offer D,16998,1,0,0,1,15,2,737.0,301.65,0.0,1010.0,1,0,92880
2257,0,0,0,0,60,1,1,DSL,0,0,1,1,One year,0,Credit card (automatic),80.55,4847.05,0,32,18,16.11,4159,0,Corona,1,0,DSL,33.833686,-117.51306299999999,0,80.55,0,0,None,21911,1,0,0,1,60,0,872.0,966.6,0.0,4847.05,0,0,92881
2258,1,0,0,0,56,1,0,DSL,1,0,0,0,One year,0,Mailed check,52.7,3019.7,0,57,27,21.61,4753,0,Corona,1,1,DSL,33.819385,-117.60021299999998,0,52.7,0,0,None,60294,0,0,0,0,56,2,0.0,1210.16,0.0,3019.7,0,1,92882
2259,0,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.85,161.65,0,31,0,11.46,4249,0,Corona,0,0,NA,33.762351,-117.488725,0,20.85,0,0,None,13188,0,0,0,0,8,0,0.0,91.68,0.0,161.65,0,0,92883
2260,0,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),80.1,217.55,1,30,64,40.67,4330,1,Yorba Linda,1,0,Cable,33.897253000000006,-117.792202,0,83.304,0,0,Offer E,39458,1,0,0,0,3,3,139.0,122.01,0.0,217.55,0,0,92886
2261,0,0,1,0,49,1,1,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),52.15,2583.75,0,19,41,28.42,5224,0,Yorba Linda,0,0,Fiber Optic,33.884073,-117.732197,1,52.15,0,6,None,20893,0,0,1,1,49,1,0.0,1392.5800000000004,0.0,2583.75,1,1,92887
2262,0,0,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.2,146.05,1,51,24,49.79,4381,1,Ventura,0,0,Cable,34.360261,-119.30638300000001,0,83.40799999999999,0,0,Offer E,32899,0,0,0,0,2,2,35.0,99.58,0.0,146.05,0,0,93001
2263,0,0,0,0,6,1,0,Fiber optic,1,1,0,1,Month-to-month,1,Bank transfer (automatic),98.15,567.45,1,20,29,20.26,3578,1,Ventura,1,0,DSL,34.279221,-119.22143700000001,0,102.076,0,0,Offer E,46894,1,0,0,1,6,2,165.0,121.56,0.0,567.45,1,0,93003
2264,1,0,0,0,70,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.95,7711.25,0,51,30,14.63,4511,0,Ventura,1,1,Fiber Optic,34.278696999999994,-119.167798,0,114.95,0,0,Offer A,27381,1,0,0,1,70,1,231.34,1024.1,0.0,7711.25,0,1,93004
2265,1,0,0,0,12,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Mailed check,112.95,1384.75,1,60,25,16.45,3965,1,Camarillo,1,1,DSL,34.227846,-119.079903,0,117.46799999999999,0,0,None,42853,1,0,0,1,12,4,346.0,197.4,0.0,1384.75,0,0,93010
2266,1,1,1,0,52,1,0,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),104.45,5481.25,0,79,11,39.0,5490,0,Camarillo,1,1,DSL,34.205504,-118.99311100000001,1,104.45,0,5,None,24945,1,0,1,0,52,0,0.0,2028.0,0.0,5481.25,0,1,93012
2267,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),113.65,8124.2,0,25,47,24.85,6469,0,Carpinteria,1,0,DSL,34.441398,-119.51316299999999,1,113.65,0,6,Offer A,17409,1,0,1,1,72,1,0.0,1789.2,0.0,8124.2,1,1,93013
2268,0,0,0,0,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.6,827.3,0,42,0,22.89,3091,0,Fillmore,0,0,NA,34.408161,-118.86511100000001,0,20.6,0,0,None,16013,0,0,0,0,40,0,0.0,915.6,0.0,827.3,0,0,93015
2269,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.9,70.9,1,43,25,39.81,4739,1,Moorpark,0,0,Cable,34.312945,-118.85816899999999,0,73.736,0,0,Offer E,32984,0,1,0,0,1,1,0.0,39.81,0.0,70.9,0,0,93021
2270,0,1,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.85,220.95,1,73,22,18.38,3561,1,Oak View,1,0,DSL,34.404544,-119.302118,0,90.324,0,0,None,6503,0,1,0,0,3,2,0.0,55.14,0.0,220.95,0,1,93022
2271,0,1,0,0,40,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,91.55,3673.6,0,72,23,44.14,5742,0,Ojai,0,0,Cable,34.581308,-118.93194799999999,0,91.55,0,0,None,21633,0,0,0,0,40,1,0.0,1765.6,0.0,3673.6,0,1,93023
2272,1,0,0,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.85,49.85,0,44,25,42.55,5323,0,Oxnard,1,1,DSL,34.223244,-119.18012,0,49.85,3,0,Offer E,79736,0,0,0,0,1,0,0.0,42.55,0.0,49.85,0,0,93030
2273,1,0,1,0,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.8,576.65,0,33,0,9.81,4006,0,Oxnard,0,1,NA,34.156628999999995,-119.117218,1,19.8,0,2,None,77791,0,0,1,0,30,2,0.0,294.3,0.0,576.65,0,0,93033
2274,1,0,1,1,23,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,99.85,2331.3,1,28,30,37.95,3425,1,Oxnard,0,1,Cable,34.184540000000005,-119.22466599999998,1,103.844,0,1,None,25322,1,0,1,1,23,1,699.0,872.85,0.0,2331.3,1,0,93035
2275,1,0,1,1,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.5,74.5,1,41,18,36.44,5554,1,Piru,0,1,DSL,34.432843,-118.730106,1,77.48,0,0,None,1459,0,1,0,0,1,2,0.0,36.44,0.0,74.5,0,1,93040
2276,0,1,1,0,44,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,104.15,4495.65,0,75,9,20.83,2944,0,Port Hueneme,1,0,DSL,34.110124,-119.100972,1,104.15,0,10,None,25634,1,0,1,0,44,1,405.0,916.52,0.0,4495.65,0,0,93041
2277,1,0,0,0,65,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,109.15,6941.2,1,60,4,9.36,6001,1,Santa Paula,1,1,Cable,34.402343,-119.094824,0,113.516,0,0,Offer B,32511,1,0,0,1,65,3,278.0,608.4,0.0,6941.2,0,0,93060
2278,0,1,0,0,7,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,48.2,340.35,0,68,21,10.53,5525,0,Simi Valley,0,0,Fiber Optic,34.296813,-118.685703,0,48.2,0,0,Offer E,49027,0,0,0,0,7,0,7.15,73.71,0.0,340.35,0,1,93063
2279,1,1,0,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.1,1789.9,0,66,0,2.37,5751,0,Simi Valley,0,1,NA,34.269449,-118.76847099999999,0,25.1,0,0,Offer A,64802,0,1,0,0,72,1,0.0,170.64,0.0,1789.9,0,0,93065
2280,0,1,0,0,8,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),100.15,908.55,0,74,23,39.86,5157,0,Somis,0,0,Fiber Optic,34.297628,-119.014627,0,100.15,0,0,Offer E,2966,1,0,0,1,8,0,20.9,318.88,0.0,908.55,0,1,93066
2281,0,0,0,0,16,1,1,DSL,0,0,0,1,Month-to-month,1,Credit card (automatic),65.2,1043.35,1,48,33,47.45,4722,1,Summerland,1,0,Cable,34.420998,-119.60136999999999,0,67.808,0,0,None,576,0,1,0,1,16,3,344.0,759.2,0.0,1043.35,0,0,93067
2282,1,1,1,1,66,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),99.5,6822.15,1,79,28,28.86,4479,1,Santa Barbara,1,1,Cable,34.419203,-119.710008,1,103.48,0,1,Offer A,31727,0,0,1,0,66,0,1910.0,1904.76,0.0,6822.15,0,0,93101
2283,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,71.55,71.55,1,42,11,17.27,5739,1,Santa Barbara,0,1,Fiber Optic,34.438581,-119.685368,0,74.41199999999999,0,0,Offer E,20893,0,0,0,0,1,0,0.0,17.27,0.0,71.55,0,0,93103
2284,1,0,0,1,3,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,55.9,157.55,0,20,69,33.28,4648,0,Santa Barbara,1,1,DSL,34.037341999999995,-119.80078999999999,0,55.9,1,0,Offer E,25771,0,0,0,1,3,1,109.0,99.84,0.0,157.55,1,0,93105
2285,1,0,1,0,53,1,1,Fiber optic,1,0,0,1,Month-to-month,0,Electronic check,93.9,5029.2,1,27,80,31.24,5543,1,Santa Barbara,1,1,DSL,34.457541,-119.631072,1,97.656,0,1,Offer B,12741,0,1,1,1,53,1,4023.0,1655.72,0.0,5029.2,1,0,93108
2286,1,1,1,0,8,1,0,DSL,0,0,0,1,Month-to-month,1,Credit card (automatic),64.4,581.7,0,78,12,25.57,4537,0,Santa Barbara,1,1,Fiber Optic,34.406256,-119.72693600000001,1,64.4,0,7,Offer E,10986,1,0,1,1,8,0,70.0,204.56,0.0,581.7,0,0,93109
2287,1,1,1,0,69,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),108.4,7318.2,1,69,4,48.88,4708,1,Santa Barbara,1,1,DSL,34.437945,-119.77191,1,112.736,0,1,Offer A,15757,1,0,1,0,69,1,293.0,3372.7200000000007,0.0,7318.2,0,0,93110
2288,0,0,0,0,5,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Mailed check,85.3,420.45,0,37,30,45.74,2689,0,Santa Barbara,0,0,DSL,34.460196999999994,-119.80260200000001,0,85.3,0,0,Offer E,16477,0,0,0,0,5,3,126.0,228.7,0.0,420.45,0,0,93111
2289,0,0,1,1,72,1,1,Fiber optic,1,0,1,1,Two year,0,Mailed check,107.45,7576.7,0,49,20,2.71,5246,0,Goleta,1,0,DSL,34.489983,-120.091246,1,107.45,2,6,Offer A,49975,1,0,1,1,72,0,1515.0,195.12,0.0,7576.7,0,0,93117
2290,0,0,1,0,13,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Bank transfer (automatic),48.75,633.4,1,42,9,0.0,2655,1,Alpaugh,1,0,Cable,35.869626000000004,-119.49877099999999,1,50.7,0,1,None,1054,0,1,1,1,13,3,0.0,0.0,0.0,633.4,0,1,93201
2291,0,0,0,0,4,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.65,321.65,1,63,22,43.32,3223,1,Armona,0,0,DSL,36.315979,-119.710852,0,89.07600000000002,0,0,Offer E,2872,0,0,0,0,4,0,71.0,173.28,0.0,321.65,0,0,93202
2292,0,0,1,1,54,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),91.3,4965,0,27,76,29.66,5907,0,Arvin,1,0,Fiber Optic,35.116307,-118.817644,1,91.3,0,5,None,16206,1,0,1,1,54,1,0.0,1601.64,0.0,4965.0,1,1,93203
2293,1,0,1,0,72,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),85.95,6151.9,0,57,30,10.97,6450,0,Avenal,1,1,DSL,35.916942999999996,-120.129921,1,85.95,0,2,Offer A,14697,1,0,1,1,72,1,0.0,789.84,0.0,6151.9,0,1,93204
2294,1,0,0,0,12,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.7,1253.9,1,44,13,25.19,2406,1,Bodfish,1,1,Cable,35.523990999999995,-118.40043200000001,0,110.96799999999999,0,0,None,1954,0,3,0,1,12,1,163.0,302.2800000000001,0.0,1253.9,0,0,93205
2295,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,25.15,25.15,1,46,6,0.0,5386,1,Buttonwillow,0,1,Cable,35.451402,-119.488413,0,26.156,0,0,Offer E,2078,0,4,0,0,1,1,0.0,0.0,0.0,25.15,0,1,93206
2296,1,1,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.2,45.2,0,73,15,49.34,4576,0,California Hot Springs,0,1,Fiber Optic,35.865795,-118.69758999999999,0,45.2,0,0,Offer E,226,0,0,0,0,1,1,0.0,49.34,0.0,45.2,0,0,93207
2297,0,0,1,0,54,1,1,Fiber optic,0,1,1,1,One year,0,Electronic check,110.35,5893.15,1,21,78,2.18,6189,1,Camp Nelson,1,0,Cable,36.057458000000004,-118.591951,1,114.764,0,1,Offer B,191,1,3,1,1,54,1,0.0,117.72,0.0,5893.15,1,1,93208
2298,1,0,1,1,69,1,1,Fiber optic,0,0,0,0,Two year,1,Credit card (automatic),79.2,5420.65,0,53,17,21.56,4072,0,Coalinga,1,1,Fiber Optic,36.186867,-120.38779299999999,1,79.2,1,5,Offer A,18036,0,0,1,0,69,0,0.0,1487.64,0.0,5420.65,0,1,93210
2299,0,0,0,0,48,1,0,DSL,1,1,0,0,Two year,0,Credit card (automatic),55.5,2627.35,0,58,5,13.03,4975,0,Corcoran,0,0,Cable,36.04533,-119.532424,0,55.5,0,0,None,23506,0,1,0,0,48,1,131.0,625.4399999999998,0.0,2627.35,0,0,93212
2300,0,0,1,1,48,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),103.25,5037.55,1,24,52,6.36,4736,1,Delano,0,0,Fiber Optic,35.772244,-119.20968899999998,1,107.38,0,1,Offer B,37280,0,0,1,1,48,4,0.0,305.2800000000001,0.0,5037.55,1,1,93215
2301,0,0,1,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,90.25,743.75,0,54,4,9.88,4969,0,Ducor,0,0,DSL,35.846067,-119.00407299999999,1,90.25,0,4,Offer E,823,1,1,1,1,8,1,30.0,79.04,0.0,743.75,0,0,93218
2302,1,0,1,1,71,1,1,DSL,1,1,1,1,Two year,1,Mailed check,91.25,6589.6,0,59,3,46.53,5529,0,Earlimart,1,1,Fiber Optic,35.858053999999996,-119.305858,1,91.25,0,7,Offer A,9318,1,1,1,1,71,2,0.0,3303.63,0.0,6589.6,0,1,93219
2303,1,0,0,0,2,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,47.8,92.45,1,35,12,13.73,4134,1,Exeter,0,1,Cable,36.301689,-119.01823300000001,0,49.712,0,0,Offer E,13333,0,0,0,0,2,1,11.0,27.46,0.0,92.45,0,0,93221
2304,1,0,1,0,67,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),100.9,6733.15,0,40,23,31.41,4078,0,Frazier Park,0,1,Fiber Optic,34.907911,-119.23428100000001,1,100.9,0,8,Offer A,1526,0,0,1,1,67,0,1549.0,2104.47,0.0,6733.15,0,0,93222
2305,1,0,1,1,34,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),97.7,3410,0,28,52,42.74,5789,0,Farmersville,0,1,Fiber Optic,36.29878,-119.20102800000001,1,97.7,2,9,None,8644,0,0,1,1,34,2,1773.0,1453.16,0.0,3410.0,1,0,93223
2306,0,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.85,199.85,0,53,21,34.76,4764,0,Fellows,0,0,Fiber Optic,35.215731,-119.57013,0,69.85,0,0,Offer E,626,0,0,0,0,3,2,42.0,104.28,0.0,199.85,0,0,93224
2307,0,0,1,1,9,1,0,DSL,0,1,1,0,One year,1,Mailed check,65.6,593.3,0,37,16,42.39,2205,0,Frazier Park,0,0,Fiber Optic,34.827662,-118.999073,1,65.6,0,2,None,4498,1,0,1,0,9,1,95.0,381.51,0.0,593.3,0,0,93225
2308,1,0,1,1,71,1,0,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),104.65,7288.4,0,23,59,14.14,6101,0,Glennville,1,1,DSL,35.735694,-118.738483,1,104.65,3,1,Offer A,296,0,0,1,1,71,2,0.0,1003.94,0.0,7288.4,1,1,93226
2309,1,0,0,0,57,1,1,Fiber optic,0,0,1,0,Two year,1,Credit card (automatic),90.45,5229.8,0,34,10,30.77,5076,0,Hanford,0,1,Fiber Optic,36.292229999999996,-119.622676,0,90.45,0,0,None,53204,1,0,0,0,57,1,523.0,1753.89,0.0,5229.8,0,0,93230
2310,1,0,0,0,72,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),63.7,4464.8,0,36,14,0.0,4921,0,Huron,1,1,Cable,36.217864,-120.08011699999999,0,63.7,0,0,Offer A,6918,1,2,0,1,72,1,0.0,0.0,0.0,4464.8,0,1,93234
2311,0,1,1,1,48,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,104.5,5068.05,0,79,75,13.4,3847,0,Ivanhoe,1,0,Fiber Optic,36.385818,-119.22424299999999,1,104.5,3,6,None,4517,1,1,1,1,48,1,0.0,643.2,0.0,5068.05,0,1,93235
2312,1,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,401.85,0,28,0,38.73,5586,0,Kernville,0,1,NA,35.852892,-118.397782,0,20.1,0,0,Offer D,1873,0,0,0,0,18,2,0.0,697.14,0.0,401.85,1,0,93238
2313,1,0,1,1,43,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),104.3,4451.85,0,20,47,22.83,3927,0,Kettleman City,1,1,Cable,35.996922999999995,-120.000951,1,104.3,2,0,None,1809,1,0,0,1,43,1,2092.0,981.69,0.0,4451.85,1,0,93239
2314,0,0,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),93.25,6688.95,0,62,7,1.72,5197,0,Lake Isabella,1,0,Fiber Optic,35.607875,-118.46631799999999,1,93.25,0,2,Offer A,5564,1,1,1,1,72,1,0.0,123.84,0.0,6688.95,0,1,93240
2315,1,0,1,1,35,1,1,DSL,0,0,1,1,One year,1,Bank transfer (automatic),73.45,2661.1,0,61,20,13.39,4719,0,Lamont,0,1,Fiber Optic,35.245034999999994,-118.905553,1,73.45,0,10,None,15364,1,0,1,1,35,0,532.0,468.65,0.0,2661.1,0,0,93241
2316,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.7,73.05,0,28,0,45.37,4676,0,Laton,0,1,NA,36.444232,-119.71828500000001,0,20.7,0,0,None,2900,0,1,0,0,4,2,0.0,181.48,0.0,73.05,1,0,93242
2317,0,0,1,1,49,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.25,1211.65,0,23,0,33.65,5616,0,Lebec,0,0,NA,34.845861,-118.88516299999999,1,25.25,2,8,None,1247,0,0,1,0,49,0,0.0,1648.85,0.0,1211.65,1,0,93243
2318,0,0,1,1,71,1,1,Fiber optic,1,1,1,0,Two year,0,Bank transfer (automatic),100.5,7030.65,0,61,19,36.5,4080,0,Lemon Cove,1,0,Cable,36.462671,-118.99729099999999,1,100.5,2,5,Offer A,293,0,1,1,0,71,3,1336.0,2591.5,0.0,7030.65,0,0,93244
2319,1,0,1,1,11,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,90.6,1020.2,0,44,19,38.48,2004,0,Lemoore,0,1,DSL,36.303666,-119.825657,1,90.6,1,9,Offer D,30419,0,0,1,1,11,1,194.0,423.28,0.0,1020.2,0,0,93245
2320,1,0,1,1,63,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),89.4,5597.65,0,39,29,44.55,5004,0,Lindsay,1,1,Fiber Optic,36.205465000000004,-119.085807,1,89.4,0,6,None,15508,1,0,1,1,63,1,1623.0,2806.65,0.0,5597.65,0,0,93247
2321,0,1,0,0,65,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),95.45,6223.3,0,69,21,32.41,4168,0,Lost Hills,1,0,Fiber Optic,35.637715,-119.893068,0,95.45,0,0,None,2502,0,2,0,0,65,1,0.0,2106.65,0.0,6223.3,0,1,93249
2322,0,0,0,1,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.45,1024.65,0,60,0,31.7,4784,0,Mc Farland,0,0,NA,35.666886,-119.18671699999999,0,20.45,3,0,None,10781,0,0,0,0,49,0,0.0,1553.3,0.0,1024.65,0,0,93250
2323,0,0,0,0,29,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),98.6,2933.2,1,49,2,27.75,5144,1,Mc Kittrick,1,0,Cable,35.38381,-119.73088500000001,0,102.544,0,0,Offer C,302,0,2,0,1,29,1,0.0,804.75,0.0,2933.2,0,1,93251
2324,0,1,1,0,15,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,83.05,1258.3,1,65,3,44.13,2596,1,Temecula,1,0,Cable,33.507255,-117.029473,1,86.37200000000001,0,2,None,46171,1,0,1,0,15,4,38.0,661.95,0.0,1258.3,0,0,92592
2325,0,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.95,82.9,0,30,0,28.55,2951,0,New Cuyama,0,0,NA,34.956577,-119.750142,1,19.95,2,1,None,798,0,0,1,0,4,2,0.0,114.2,0.0,82.9,0,0,93254
2326,0,0,1,0,72,1,1,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),109.15,7789.6,0,21,82,11.85,4807,0,Temecula,1,0,Fiber Optic,33.507255,-117.029473,1,109.15,0,2,Offer A,46171,1,0,1,1,72,0,0.0,853.1999999999998,0.0,7789.6,1,1,92592
2327,0,1,1,0,26,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),85.7,2067,0,68,4,46.24,3935,0,Pixley,1,0,Fiber Optic,35.957019,-119.330928,1,85.7,0,4,None,4198,0,0,1,0,26,0,0.0,1202.24,0.0,2067.0,0,1,93256
2328,0,1,1,0,35,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),102.05,3452.55,0,70,10,45.13,3199,0,Porterville,1,0,Cable,36.008958,-118.891593,1,102.05,0,1,None,65566,0,0,1,1,35,0,345.0,1579.5500000000004,0.0,3452.55,0,0,93257
2329,0,0,0,0,57,1,1,Fiber optic,0,1,0,1,One year,0,Electronic check,94.7,5468.95,0,47,7,38.94,4507,0,Posey,0,0,Cable,35.861928000000006,-118.636698,0,94.7,0,0,None,266,1,0,0,1,57,0,383.0,2219.58,0.0,5468.95,0,0,93260
2330,1,0,1,1,28,1,1,DSL,0,1,0,1,Month-to-month,0,Electronic check,64.4,1802.15,0,52,19,9.31,2434,0,Richgrove,0,1,DSL,35.809921,-119.12743700000001,1,64.4,2,2,None,2956,0,0,1,1,28,1,342.0,260.68,0.0,1802.15,0,0,93261
2331,0,0,1,0,25,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,26.8,733.55,0,56,0,3.6,3428,0,Sequoia National Park,0,0,NA,36.527243,-118.59493799999998,1,26.8,0,10,None,56,0,0,1,0,25,2,0.0,90.0,0.0,733.55,0,0,93262
2332,0,0,1,0,47,1,0,DSL,1,0,1,0,One year,1,Credit card (automatic),66.05,3021.45,0,49,11,6.56,3404,0,Shafter,1,0,Fiber Optic,35.490705,-119.286833,1,66.05,0,1,None,15177,0,0,1,0,47,0,0.0,308.32,0.0,3021.45,0,1,93263
2333,0,0,1,1,57,1,1,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),65.2,3687.85,0,35,15,1.54,4491,0,Springville,0,0,Fiber Optic,36.245926000000004,-118.69313799999999,1,65.2,1,3,None,3546,1,0,1,0,57,1,0.0,87.78,0.0,3687.85,0,1,93265
2334,1,1,1,0,16,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),85.05,1391.15,0,69,6,48.41,3739,0,Stratford,0,1,DSL,36.175255,-119.813805,1,85.05,0,6,Offer D,1729,0,0,1,0,16,0,83.0,774.56,0.0,1391.15,0,0,93266
2335,1,0,0,0,5,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,55.8,274.35,0,24,51,41.29,2612,0,Strathmore,1,1,Cable,36.141319,-119.129075,0,55.8,0,0,None,5689,0,1,0,0,5,1,140.0,206.45,0.0,274.35,1,0,93267
2336,1,0,1,0,17,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),70.4,1214.05,1,35,12,13.68,4469,1,Taft,0,1,Fiber Optic,35.184837,-119.402525,1,73.21600000000002,0,1,None,14937,0,1,1,0,17,3,146.0,232.56,0.0,1214.05,0,0,93268
2337,0,1,0,0,56,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),104.75,5510.65,1,68,4,34.58,5605,1,Terra Bella,1,0,DSL,35.939068,-119.04366599999999,0,108.94,0,0,None,5868,0,0,0,0,56,2,0.0,1936.48,0.0,5510.65,0,1,93270
2338,1,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.95,1322.85,0,48,0,8.53,5092,0,Three Rivers,0,1,NA,36.413433000000005,-118.854708,1,19.95,2,0,Offer A,2318,0,2,0,0,72,2,0.0,614.16,0.0,1322.85,0,0,93271
2339,0,1,0,0,21,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.25,1973.75,1,79,10,21.15,4819,1,Temecula,0,0,DSL,33.507255,-117.029473,0,98.02,0,0,None,46171,0,0,0,0,21,0,197.0,444.15,0.0,1973.75,0,0,92592
2340,0,0,1,1,48,0,No phone service,DSL,1,0,0,1,One year,0,Credit card (automatic),45.0,2196.3,0,43,22,0.0,5269,0,Tulare,1,0,Fiber Optic,36.185471,-119.375243,1,45.0,3,3,None,56101,0,0,1,1,48,3,0.0,0.0,0.0,2196.3,0,1,93274
2341,0,0,1,0,68,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),114.9,7843.55,0,46,21,23.14,5782,0,Tupman,1,0,Fiber Optic,35.316263,-119.40255900000001,1,114.9,0,8,Offer A,236,1,0,1,1,68,2,1647.0,1573.52,0.0,7843.55,0,0,93276
2342,0,0,0,0,30,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Bank transfer (automatic),106.4,3211.9,0,22,73,42.49,5503,0,Visalia,0,0,Fiber Optic,36.303793,-119.375646,0,106.4,0,0,None,44741,1,0,0,1,30,0,2345.0,1274.7,0.0,3211.9,1,0,93277
2343,0,0,1,0,3,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,46.1,130.15,0,61,7,2.66,4047,0,Wasco,0,0,DSL,35.652242,-119.4464,1,46.1,0,2,None,22760,0,0,1,0,3,0,0.0,7.98,0.0,130.15,0,1,93280
2344,0,1,0,0,14,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,39.7,692.35,0,75,24,0.0,3162,0,Weldon,1,0,Fiber Optic,35.556470000000004,-118.244914,0,39.7,0,0,Offer D,1935,1,0,0,0,14,2,166.0,0.0,0.0,692.35,0,0,93283
2345,0,0,0,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.05,85.5,0,57,0,27.37,4462,0,Wofford Heights,0,0,NA,35.690535,-118.552784,0,20.05,2,0,None,2515,0,0,0,0,4,0,0.0,109.48,0.0,85.5,0,0,93285
2346,0,0,1,1,71,1,1,Fiber optic,0,1,0,1,Two year,1,Credit card (automatic),95.75,6849.4,0,58,12,27.26,4865,0,Woodlake,1,0,Fiber Optic,36.464634999999994,-119.094348,1,95.75,2,9,Offer A,8870,0,0,1,1,71,2,822.0,1935.46,0.0,6849.4,0,0,93286
2347,1,0,1,1,8,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,24.4,203.95,0,43,0,23.18,2028,0,Woody,0,1,NA,35.710244,-118.881679,1,24.4,0,6,None,88,0,0,1,0,8,1,0.0,185.44,0.0,203.95,0,0,93287
2348,1,0,1,1,61,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),33.6,2117.2,0,24,76,0.0,6495,0,Visalia,1,1,DSL,36.391777000000005,-119.37284199999999,1,33.6,1,3,None,36718,0,0,1,0,61,0,0.0,0.0,0.0,2117.2,1,1,93291
2349,1,0,1,1,72,1,1,Fiber optic,0,1,0,0,Two year,0,Bank transfer (automatic),90.45,6565.85,0,31,24,8.51,4461,0,Visalia,1,1,Fiber Optic,36.37559,-119.21168899999999,1,90.45,3,7,Offer A,30395,1,0,1,0,72,1,1576.0,612.72,0.0,6565.85,0,0,93292
2350,0,0,0,0,5,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.0,424.75,0,29,85,48.49,4456,0,Bakersfield,0,0,Fiber Optic,35.383937,-119.02042800000001,0,84.0,0,0,None,12963,0,0,0,0,5,1,361.0,242.45,0.0,424.75,1,0,93301
2351,0,0,0,0,49,1,0,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),67.4,3306.85,0,37,23,20.45,5075,0,Bakersfield,1,0,Cable,35.339796,-119.023552,0,67.4,0,0,None,44588,1,0,0,0,49,2,0.0,1002.05,0.0,3306.85,0,1,93304
2352,1,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.7,168.9,0,28,0,22.15,5498,0,Bakersfield,0,1,NA,35.391733,-118.984109,0,19.7,0,0,Offer E,35643,0,0,0,0,8,1,0.0,177.2,0.0,168.9,1,0,93305
2353,1,0,0,0,3,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.35,253.8,0,60,26,49.63,4203,0,Bakersfield,0,1,DSL,35.449881,-118.84144199999999,0,80.35,0,0,Offer E,53481,0,0,0,1,3,0,66.0,148.89,0.0,253.8,0,0,93306
2354,1,0,1,1,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.6,197.4,0,53,0,2.68,4406,0,Bakersfield,0,1,NA,35.280113,-118.962329,1,19.6,3,9,Offer E,59195,0,0,1,0,9,0,0.0,24.12,0.0,197.4,0,0,93307
2355,1,0,1,1,67,1,0,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),54.2,3838.2,0,42,26,10.9,6005,0,Bakersfield,0,1,DSL,35.559616999999996,-118.92518500000001,1,54.2,2,1,Offer A,44915,0,0,1,0,67,0,0.0,730.3000000000002,0.0,3838.2,0,1,93308
2356,1,0,0,0,46,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),45.2,2065.15,0,36,16,24.13,3150,0,Bakersfield,0,1,Fiber Optic,35.342890999999995,-119.064803,0,45.2,0,0,Offer B,58632,0,0,0,0,46,1,330.0,1109.98,0.0,2065.15,0,0,93309
2357,0,0,1,0,67,1,1,DSL,1,1,0,1,One year,0,Mailed check,75.1,5064.45,0,23,58,4.71,4931,0,Bakersfield,1,0,Cable,35.16207,-119.19448799999999,1,75.1,0,10,Offer A,20440,0,0,1,1,67,1,2937.0,315.57,0.0,5064.45,1,0,93311
2358,0,0,1,0,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.7,1140.05,0,54,0,3.28,4888,0,Bakersfield,0,0,NA,35.392599,-119.245341,1,19.7,0,8,Offer B,40836,0,0,1,0,55,0,0.0,180.4,0.0,1140.05,0,0,93312
2359,1,0,1,0,33,1,1,DSL,1,1,1,0,Month-to-month,1,Bank transfer (automatic),72.75,2447.45,0,54,21,19.11,4959,0,Bakersfield,1,1,Fiber Optic,35.140938,-119.051348,1,72.75,0,1,None,25126,0,0,1,0,33,1,51.4,630.63,0.0,2447.45,0,1,93313
2360,1,0,1,1,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.05,1263.9,0,64,0,20.96,6444,0,San Luis Obispo,0,1,NA,35.233745,-120.626442,1,20.05,1,5,Offer B,27047,0,0,1,0,62,0,0.0,1299.52,0.0,1263.9,0,0,93401
2361,0,0,0,1,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.95,45.95,1,49,21,46.17,4563,1,Los Osos,0,0,Cable,35.279984000000006,-120.824288,0,47.788,1,0,Offer E,14859,0,2,0,0,1,1,0.0,46.17,0.0,45.95,0,0,93402
2362,1,0,1,1,49,0,No phone service,DSL,1,0,0,1,Month-to-month,1,Electronic check,39.2,1838.15,0,24,47,0.0,4810,0,San Luis Obispo,0,1,Cable,35.236549,-120.72734399999999,1,39.2,2,8,Offer B,31982,0,0,1,1,49,0,864.0,0.0,0.0,1838.15,1,0,93405
2363,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.75,44.75,0,37,26,18.57,5479,0,Arroyo Grande,0,1,Fiber Optic,35.176235999999996,-120.48324299999999,0,44.75,0,0,Offer E,24499,0,0,0,0,1,2,0.0,18.57,0.0,44.75,0,0,93420
2364,1,0,1,0,14,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,82.65,1185,0,37,10,45.57,4965,0,Atascadero,1,1,DSL,35.453912,-120.69461000000001,1,82.65,0,8,Offer D,29539,0,0,1,0,14,2,118.0,637.98,0.0,1185.0,0,0,93422
2365,1,1,0,0,18,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Bank transfer (automatic),93.9,1743.9,0,75,25,1.92,3728,0,Avila Beach,1,1,DSL,35.186644,-120.728305,0,93.9,0,0,Offer D,812,1,0,0,0,18,1,436.0,34.56,0.0,1743.9,0,0,93424
2366,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.15,70.15,1,80,9,47.97,2825,1,Bradley,0,0,Fiber Optic,35.842889,-121.00486200000002,0,72.956,0,0,None,1363,0,0,0,0,1,1,0.0,47.97,0.0,70.15,0,1,93426
2367,0,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),85.55,85.55,1,45,4,33.34,3967,1,Buellton,1,0,DSL,34.631362,-120.23821799999999,0,88.97200000000001,0,0,Offer E,4644,0,0,0,0,1,1,0.0,33.34,0.0,85.55,0,0,93427
2368,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),117.15,8529.5,0,43,5,24.89,4743,0,Cambria,1,0,Cable,35.591387,-121.032256,1,117.15,0,1,Offer A,6526,1,0,1,1,72,2,42.65,1792.08,0.0,8529.5,0,1,93428
2369,1,0,0,0,64,1,1,Fiber optic,1,0,0,1,Two year,0,Credit card (automatic),99.25,6549.45,0,38,14,36.54,5213,0,Casmalia,1,1,DSL,34.866032000000004,-120.536546,0,99.25,0,0,Offer B,210,1,0,0,1,64,0,91.69,2338.56,0.0,6549.45,0,1,93429
2370,1,0,1,0,69,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),112.55,7806.5,0,29,41,3.41,5532,0,Cayucos,1,1,Fiber Optic,35.511833,-120.91871299999998,1,112.55,0,9,Offer A,3220,1,0,1,1,69,0,0.0,235.29,0.0,7806.5,1,1,93430
2371,0,0,0,0,1,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,25.7,25.7,0,30,0,43.84,5249,0,Creston,0,0,NA,35.480896,-120.469476,0,25.7,0,0,Offer E,1203,0,0,0,0,1,0,0.0,43.84,0.0,25.7,0,0,93432
2372,1,0,1,1,71,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),90.3,6287.3,0,48,57,15.71,6291,0,Grover Beach,1,1,Cable,35.120833000000005,-120.61843,1,90.3,3,1,Offer A,13106,1,1,1,1,71,1,3584.0,1115.41,0.0,6287.3,0,0,93433
2373,0,0,1,1,66,1,0,DSL,0,0,0,0,One year,1,Credit card (automatic),49.4,3251.85,0,34,27,48.11,5232,0,Guadalupe,0,0,Cable,34.936,-120.594655,1,49.4,2,1,Offer A,5726,1,0,1,0,66,0,0.0,3175.26,0.0,3251.85,0,1,93434
2374,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.4,50.6,0,32,0,15.16,3954,0,Lompoc,0,1,NA,34.601055,-120.38291699999999,0,19.4,0,0,Offer E,51737,0,0,0,0,2,0,0.0,30.32,0.0,50.6,0,0,93436
2375,0,1,1,0,71,1,0,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),109.7,7904.25,0,67,14,9.96,5011,0,Lompoc,1,0,Fiber Optic,34.757477,-120.55050700000001,1,109.7,0,1,Offer A,6165,1,0,1,1,71,0,0.0,707.1600000000002,0.0,7904.25,0,1,93437
2376,1,0,0,0,11,1,0,DSL,0,1,1,0,One year,1,Electronic check,61.25,729.95,0,29,59,27.84,2738,0,Los Alamos,0,1,Cable,34.758699,-120.27583899999999,0,61.25,0,0,Offer D,1328,0,0,0,0,11,0,431.0,306.24,0.0,729.95,1,0,93440
2377,1,0,0,1,47,1,0,DSL,1,1,0,0,Month-to-month,1,Electronic check,55.3,2654.05,0,52,17,25.25,5491,0,Los Olivos,0,1,Cable,34.70434,-120.02609,0,55.3,2,0,Offer B,1317,0,0,0,0,47,0,0.0,1186.75,0.0,2654.05,0,1,93441
2378,0,0,1,0,35,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,2416.55,1,61,4,10.43,5413,1,Morro Bay,0,0,Fiber Optic,35.369553,-120.76386399999998,1,73.112,0,4,Offer C,10909,0,0,1,0,35,1,97.0,365.05,0.0,2416.55,0,0,93442
2379,1,1,1,0,32,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Bank transfer (automatic),106.35,3520.75,1,77,3,7.92,4113,1,Nipomo,1,1,Cable,35.050345,-120.489599,1,110.604,0,3,None,15405,0,1,1,0,32,3,106.0,253.44,0.0,3520.75,0,0,93444
2380,1,0,1,1,60,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),103.75,5969.95,0,57,19,2.83,6237,0,Oceano,0,1,Fiber Optic,35.059695,-120.60474099999999,1,103.75,1,1,Offer B,7435,1,1,1,1,60,2,1134.0,169.8,0.0,5969.95,0,0,93445
2381,1,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.5,226.8,0,22,0,33.48,5825,0,Paso Robles,0,1,NA,35.634221999999994,-120.72834099999999,0,19.5,0,0,Offer D,35586,0,0,0,0,11,1,0.0,368.28,0.0,226.8,1,0,93446
2382,0,0,0,0,29,0,No phone service,DSL,1,1,0,0,One year,0,Credit card (automatic),39.5,1082.75,0,47,28,0.0,5103,0,Pismo Beach,0,0,DSL,35.165668,-120.65584199999999,0,39.5,0,0,None,8564,1,0,0,0,29,2,0.0,0.0,0.0,1082.75,0,1,93449
2383,1,0,1,1,21,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,26.05,565.75,0,23,59,0.0,4302,0,San Ardo,0,1,DSL,35.996008,-120.85305,1,26.05,9,1,Offer D,670,0,0,1,0,21,2,334.0,0.0,0.0,565.75,1,0,93450
2384,1,1,1,0,48,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),91.05,4370.75,0,65,22,25.19,3594,0,San Miguel,1,1,DSL,35.886767,-120.60866100000001,1,91.05,0,1,None,2666,0,0,1,1,48,0,0.0,1209.12,0.0,4370.75,0,1,93451
2385,0,0,0,1,3,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Mailed check,29.65,90.05,0,44,53,0.0,5880,0,San Simeon,0,0,Fiber Optic,35.746484,-121.223355,0,29.65,3,0,None,471,0,0,0,0,3,0,0.0,0.0,0.0,90.05,0,1,93452
2386,0,0,1,1,43,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,50.2,2169.4,0,41,19,14.64,5284,0,Santa Margarita,0,0,DSL,35.303926000000004,-120.25656699999999,1,50.2,2,1,Offer B,2687,0,0,1,0,43,0,412.0,629.52,0.0,2169.4,0,0,93453
2387,1,0,0,0,5,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,105.3,550.6,0,34,30,44.65,4024,0,Santa Maria,1,1,DSL,34.943523,-120.256729,0,105.3,0,0,Offer E,30540,0,0,0,1,5,0,0.0,223.25,0.0,550.6,0,1,93454
2388,0,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.45,55.45,0,63,27,6.43,5286,0,Santa Maria,0,0,Fiber Optic,34.818227,-120.418784,0,55.45,0,0,Offer E,37364,0,0,0,1,1,2,0.0,6.43,0.0,55.45,0,1,93455
2389,1,0,1,1,71,1,1,DSL,1,0,1,1,One year,0,Electronic check,85.45,6300.85,0,57,53,23.41,5280,0,Santa Maria,1,1,DSL,34.959340000000005,-120.490081,1,85.45,3,0,Offer A,43684,1,1,0,1,71,1,0.0,1662.11,0.0,6300.85,0,1,93458
2390,0,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.8,160.05,0,20,0,28.37,5698,0,Santa Ynez,0,0,NA,34.630356,-120.032564,1,19.8,0,1,Offer E,5710,0,0,1,0,8,2,0.0,226.96,0.0,160.05,1,0,93460
2391,1,0,0,0,8,1,1,DSL,0,0,1,0,Month-to-month,1,Electronic check,59.25,436.6,0,38,22,48.2,3003,0,Shandon,0,1,Cable,35.634488,-120.29353400000001,0,59.25,0,0,Offer E,1255,0,0,0,0,8,1,0.0,385.6,0.0,436.6,0,1,93461
2392,1,0,0,0,20,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),90.7,1781.35,0,38,27,25.41,2927,0,Solvang,1,1,Cable,34.624399,-120.137875,0,90.7,0,0,Offer D,7958,0,1,0,0,20,4,481.0,508.2,0.0,1781.35,0,0,93463
2393,0,0,1,1,33,1,1,Fiber optic,1,0,1,1,One year,1,Mailed check,103.7,3467,1,22,80,41.61,4461,1,Templeton,1,0,DSL,35.536115,-120.739231,1,107.848,0,1,Offer C,7918,0,2,1,1,33,2,2774.0,1373.13,0.0,3467.0,1,0,93465
2394,1,0,0,0,71,1,1,Fiber optic,0,1,0,0,One year,1,Credit card (automatic),79.05,5552.5,0,44,10,41.34,5466,0,Mojave,0,1,Fiber Optic,35.097322999999996,-118.17128799999999,0,79.05,0,0,Offer A,4882,0,0,0,0,71,0,0.0,2935.140000000001,0.0,5552.5,0,1,93501
2395,0,1,1,0,31,1,1,Fiber optic,0,0,1,0,One year,1,Electronic check,90.7,2835.5,0,67,22,44.26,2364,0,California City,1,0,DSL,35.151491,-117.92759699999999,1,90.7,0,1,None,8316,0,0,1,0,31,0,0.0,1372.06,0.0,2835.5,0,1,93505
2396,0,1,1,0,38,1,1,Fiber optic,1,1,0,1,One year,0,Credit card (automatic),95.0,3591.25,0,74,27,49.82,5148,0,Acton,0,0,DSL,34.501452,-118.207862,1,95.0,0,1,None,7831,0,0,1,1,38,0,970.0,1893.16,0.0,3591.25,0,0,93510
2397,1,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,88.35,88.35,1,23,51,14.26,4254,1,Benton,0,1,Cable,37.653946999999995,-118.231443,0,91.884,0,0,None,340,0,0,0,1,1,3,0.0,14.26,0.0,88.35,1,0,93512
2398,0,0,1,1,2,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Mailed check,30.25,63.75,0,31,20,0.0,4387,0,Big Pine,0,0,Fiber Optic,37.245505,-118.06294299999999,1,30.25,2,6,Offer E,1826,0,2,1,0,2,3,0.0,0.0,0.0,63.75,0,1,93513
2399,0,0,1,0,12,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Bank transfer (automatic),49.85,617.15,0,24,82,0.0,2873,0,Bishop,1,0,Fiber Optic,37.045840000000005,-118.397236,1,49.85,0,10,Offer D,13309,0,0,1,1,12,0,0.0,0.0,0.0,617.15,1,1,93514
2400,0,0,0,1,9,1,0,Fiber optic,1,0,0,1,Month-to-month,0,Bank transfer (automatic),93.0,870.25,0,46,16,42.1,2267,0,Boron,1,0,Fiber Optic,34.957029999999996,-117.73045,0,93.0,1,0,None,2241,1,0,0,1,9,2,139.0,378.9,0.0,870.25,0,0,93516
2401,1,1,0,1,11,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,54.55,601.25,0,72,23,11.86,4143,0,Bridgeport,0,1,Fiber Optic,38.184583,-119.28655800000001,0,54.55,1,0,None,826,1,0,0,0,11,0,0.0,130.45999999999998,0.0,601.25,0,1,93517
2402,1,0,0,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.7,111.65,0,46,0,27.78,2276,0,Caliente,0,1,NA,35.358953,-118.527064,0,19.7,1,0,None,1022,0,0,0,0,6,3,0.0,166.68,0.0,111.65,0,0,93518
2403,0,0,1,0,71,1,0,DSL,1,1,1,1,One year,1,Bank transfer (automatic),84.8,6046.1,0,50,6,23.06,5643,0,Darwin,1,0,DSL,36.319181,-117.593053,1,84.8,0,2,None,64,1,0,1,1,71,0,36.28,1637.26,0.0,6046.1,0,1,93522
2404,0,0,1,1,42,1,1,Fiber optic,1,1,1,0,One year,1,Credit card (automatic),94.45,3923.8,0,21,69,6.37,5643,0,Edwards,0,0,DSL,34.966777,-117.961179,1,94.45,3,5,Offer B,7685,0,0,1,0,42,0,2707.0,267.54,0.0,3923.8,1,0,93523
2405,0,0,1,1,8,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.2,777.3,1,22,84,38.83,2939,1,Independence,1,0,Fiber Optic,36.869584,-118.189241,1,97.96799999999999,0,1,Offer E,734,0,3,1,1,8,1,653.0,310.64,0.0,777.3,1,0,93526
2406,0,0,0,0,5,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,96.25,512.45,1,62,11,32.12,5056,1,Temecula,0,0,Cable,33.507255,-117.029473,0,100.1,0,0,Offer E,46171,0,0,0,1,5,4,56.0,160.6,0.0,512.45,0,0,92592
2407,0,0,1,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.7,141.45,1,28,30,9.76,4559,1,San Diego,0,0,Fiber Optic,32.961064,-117.13491699999999,1,73.528,0,1,Offer E,47224,0,0,1,0,2,4,42.0,19.52,0.0,141.45,1,0,92129
2408,0,0,1,1,45,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.85,892.15,0,24,0,40.19,2844,0,June Lake,0,0,NA,37.730269,-119.05581299999999,1,20.85,1,2,Offer B,618,0,0,1,0,45,1,0.0,1808.55,0.0,892.15,1,0,93529
2409,1,0,1,1,28,0,No phone service,DSL,0,1,1,1,One year,1,Credit card (automatic),60.0,1682.05,0,58,52,0.0,2797,0,Keeler,1,1,Cable,36.560497999999995,-117.962461,1,60.0,3,8,None,71,1,1,1,1,28,2,875.0,0.0,0.0,1682.05,0,0,93530
2410,0,0,1,0,43,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,80.45,3398.9,0,41,15,41.83,5357,0,Keene,0,0,Fiber Optic,35.214982,-118.59048999999999,1,80.45,0,7,Offer B,1436,0,0,1,0,43,1,510.0,1798.6899999999996,0.0,3398.9,0,0,93531
2411,1,0,0,1,60,1,1,DSL,1,0,1,1,Two year,1,Electronic check,84.95,4984.85,0,28,85,49.96,4104,0,Lake Hughes,1,1,Cable,34.659579,-118.58421200000001,0,84.95,1,0,Offer B,2771,1,0,0,1,60,0,423.71,2997.6,0.0,4984.85,1,1,93532
2412,0,0,1,0,42,0,No phone service,DSL,0,1,0,0,One year,0,Mailed check,33.55,1445.3,1,55,6,0.0,2044,1,Lancaster,0,0,Fiber Optic,34.727529,-118.153098,1,34.892,0,1,Offer B,35109,1,1,1,0,42,1,87.0,0.0,0.0,1445.3,0,0,93534
2413,1,0,1,1,7,0,No phone service,DSL,1,0,0,1,Two year,0,Credit card (automatic),49.65,305.55,0,46,28,0.0,2750,0,Lancaster,1,1,Fiber Optic,34.712708,-117.889656,1,49.65,2,4,None,57794,1,0,1,1,7,1,86.0,0.0,0.0,305.55,0,0,93535
2414,0,0,1,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.2,507.9,0,21,0,10.49,4129,0,Lancaster,0,0,NA,34.741406,-118.38111,1,20.2,0,2,None,49309,0,0,1,0,25,1,0.0,262.25,0.0,507.9,1,0,93536
2415,0,1,1,1,40,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),94.55,3640.45,1,65,22,49.5,5676,1,Lee Vining,0,0,Cable,37.890145000000004,-119.184087,1,98.33200000000001,0,1,None,504,0,2,1,1,40,3,0.0,1980.0,0.0,3640.45,0,1,93541
2416,1,0,0,0,27,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),100.5,2673.45,0,23,73,8.86,5939,0,Littlerock,1,1,DSL,34.505272999999995,-117.955054,0,100.5,0,0,Offer C,11198,0,0,0,1,27,0,0.0,239.22,0.0,2673.45,1,1,93543
2417,1,0,0,0,10,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,35.75,389.8,0,53,22,0.0,2263,0,Llano,0,1,Cable,34.500091,-117.76586200000001,0,35.75,0,0,Offer D,1220,1,0,0,0,10,4,0.0,0.0,0.0,389.8,0,1,93544
2418,0,1,0,0,27,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),86.45,2401.05,0,77,4,2.97,5990,0,Fallbrook,1,0,Cable,33.362575,-117.299644,0,86.45,0,0,None,42239,0,0,0,0,27,1,96.0,80.19000000000003,0.0,2401.05,0,0,92028
2419,0,0,0,0,11,1,0,DSL,0,0,0,0,One year,0,Bank transfer (automatic),53.8,651.55,0,33,17,7.42,5899,0,Mammoth Lakes,1,0,DSL,37.550074,-118.837167,0,53.8,0,0,Offer D,8217,1,0,0,0,11,2,111.0,81.62,0.0,651.55,0,0,93546
2420,1,0,1,1,4,0,No phone service,DSL,1,0,1,0,Month-to-month,0,Credit card (automatic),38.55,156.1,0,56,53,0.0,3824,0,Olancha,0,1,Cable,36.296851000000004,-117.86546899999999,1,38.55,3,3,None,318,0,0,1,0,4,0,83.0,0.0,0.0,156.1,0,0,93549
2421,1,0,0,0,68,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Bank transfer (automatic),39.9,2796.35,0,19,58,0.0,6270,0,Palmdale,1,1,DSL,34.536232,-118.082935,0,39.9,0,0,None,67232,0,0,0,1,68,3,1622.0,0.0,0.0,2796.35,1,0,93550
2422,1,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.05,70.05,0,72,5,2.97,2469,0,Palmdale,0,1,DSL,34.613476,-118.256358,0,70.05,0,0,Offer E,34045,0,0,0,0,1,0,0.0,2.97,0.0,70.05,0,0,93551
2423,0,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,407.05,0,38,0,18.8,2910,0,Palmdale,0,0,NA,34.557711,-118.02944099999999,0,20.1,0,0,Offer D,25370,0,0,0,0,18,1,0.0,338.4000000000001,0.0,407.05,0,0,93552
2424,0,0,0,0,57,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),112.95,6465,1,38,7,48.86,4738,1,Pearblossom,1,0,Cable,34.445239,-117.89486799999999,0,117.46799999999999,0,0,None,1613,0,0,0,1,57,1,0.0,2785.02,0.0,6465.0,0,1,93553
2425,1,0,0,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.3,511.25,0,57,0,13.34,5712,0,Randsburg,0,1,NA,35.405722,-117.773354,0,20.3,0,0,Offer C,117,0,0,0,0,26,2,0.0,346.84,0.0,511.25,0,0,93554
2426,0,0,1,0,17,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),35.65,646.05,0,48,23,0.0,5977,0,Temecula,1,0,Fiber Optic,33.507255,-117.029473,1,35.65,0,5,Offer D,46171,0,0,1,0,17,1,0.0,0.0,0.0,646.05,0,1,92592
2427,1,0,0,0,1,0,No phone service,DSL,0,0,0,1,Month-to-month,0,Electronic check,35.9,35.9,1,54,32,0.0,4747,1,Rosamond,0,1,Cable,34.903052,-118.41125100000001,0,37.336,0,0,Offer E,14931,0,4,0,1,1,4,0.0,0.0,0.0,35.9,0,1,93560
2428,1,0,0,1,38,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),99.25,3777.15,1,30,94,31.27,5274,1,Tehachapi,1,1,Fiber Optic,35.073777,-118.65211200000002,0,103.22,0,0,Offer C,25805,0,2,0,1,38,4,355.05,1188.26,0.0,3777.15,0,1,93561
2429,1,1,1,0,59,1,0,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),82.95,4903.15,0,75,21,4.21,5295,0,Temecula,1,1,Cable,33.507255,-117.029473,1,82.95,0,10,None,46171,0,0,1,0,59,0,1030.0,248.39,0.0,4903.15,0,0,92592
2430,1,0,0,0,30,1,0,DSL,1,0,0,0,Two year,1,Mailed check,55.65,1653.85,0,35,24,47.06,5445,0,Valyermo,1,1,Fiber Optic,34.39583,-117.734568,0,55.65,0,0,Offer C,413,0,0,0,0,30,0,39.69,1411.8000000000004,0.0,1653.85,0,1,93563
2431,1,1,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,24.45,47.5,1,66,7,0.0,5573,1,Palmdale,0,1,DSL,34.598221,-117.79593,0,25.428,0,0,None,6787,0,0,0,0,2,3,3.0,0.0,0.0,47.5,0,0,93591
2432,0,1,1,0,50,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,25.2,1306.3,0,79,0,31.43,4015,0,Ahwahnee,0,0,NA,37.375816,-119.739935,1,25.2,0,0,None,1968,0,0,0,0,50,4,0.0,1571.5,0.0,1306.3,0,0,93601
2433,1,0,0,0,9,0,No phone service,DSL,1,0,0,1,One year,0,Mailed check,50.8,463.6,0,61,14,0.0,5535,0,Auberry,1,1,Fiber Optic,36.991762,-119.242874,0,50.8,0,0,None,3464,1,0,0,1,9,2,65.0,0.0,0.0,463.6,0,0,93602
2434,0,0,1,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,60.65,0,44,0,30.34,4943,0,Badger,0,0,NA,36.64545,-118.924982,1,19.65,3,1,None,273,0,0,1,0,3,0,0.0,91.02,0.0,60.65,0,0,93603
2435,0,0,0,1,14,1,0,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),59.8,824.85,0,44,24,44.14,5962,0,Bass Lake,1,0,DSL,37.458366999999996,-119.34501100000001,0,59.8,1,0,Offer D,613,0,0,0,0,14,0,19.8,617.96,0.0,824.85,0,1,93604
2436,0,1,0,0,31,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),73.55,2094.65,0,72,8,47.48,2057,0,Big Creek,0,0,Fiber Optic,37.17277,-119.2997,0,73.55,0,0,None,273,0,0,0,0,31,3,168.0,1471.88,0.0,2094.65,0,0,93605
2437,0,0,0,0,7,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,61.4,438.9,0,38,14,15.84,2845,0,Biola,1,0,Fiber Optic,36.798882,-120.01951100000001,0,61.4,0,0,None,807,0,0,0,0,7,0,0.0,110.88,0.0,438.9,0,1,93606
2438,0,0,0,0,8,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),103.35,847.3,1,26,45,19.68,2363,1,Cantua Creek,0,0,DSL,36.488056,-120.40769099999999,0,107.484,0,0,Offer E,1766,1,0,0,1,8,2,381.0,157.44,0.0,847.3,1,0,93608
2439,1,0,1,1,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.9,329.75,0,61,0,14.69,3526,0,Caruthers,0,1,NA,36.5276,-119.865999,1,19.9,0,8,Offer D,5446,0,0,1,0,17,1,0.0,249.73,0.0,329.75,0,0,93609
2440,1,0,1,1,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.45,674.55,0,22,0,35.05,4363,0,Chowchilla,0,1,NA,37.100947999999995,-120.27013600000001,1,19.45,3,5,Offer C,19391,0,0,1,0,32,0,0.0,1121.6,0.0,674.55,1,0,93610
2441,0,1,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Mailed check,81.5,162.55,0,66,22,24.95,4267,0,Clovis,0,0,DSL,36.917652000000004,-119.59375700000001,0,81.5,0,0,None,46858,0,0,0,0,2,0,36.0,49.9,0.0,162.55,0,0,93611
2442,1,1,0,0,7,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.8,546.95,1,75,14,39.51,2015,1,Clovis,0,1,Cable,36.814539,-119.711868,0,88.19200000000001,0,0,None,33856,0,0,0,0,7,6,0.0,276.57,0.0,546.95,0,1,93612
2443,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),109.55,7887.25,0,27,52,33.39,5723,0,Coarsegold,1,0,Cable,37.212191,-119.749323,1,109.55,3,9,None,9395,0,0,1,1,72,0,4101.0,2404.08,0.0,7887.25,1,0,93614
2444,0,1,0,0,31,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.95,3186.65,1,74,4,39.36,5362,1,Cutler,0,0,Fiber Optic,36.497895,-119.28548400000001,0,103.948,0,0,None,5519,0,0,0,0,31,4,12.75,1220.16,0.0,3186.65,0,1,93615
2445,0,0,1,1,27,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Mailed check,74.4,1972.35,0,56,28,46.66,4331,0,Del Rey,0,0,Fiber Optic,36.657462,-119.595293,1,74.4,2,6,Offer C,1965,0,0,1,0,27,1,0.0,1259.82,0.0,1972.35,0,1,93616
2446,0,0,0,0,18,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),90.0,1527.35,1,55,6,13.65,2708,1,Dinuba,0,0,Cable,36.523619000000004,-119.38686799999999,0,93.6,0,0,None,24206,0,0,0,0,18,0,0.0,245.7,0.0,1527.35,0,1,93618
2447,1,0,0,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.9,490.55,0,55,12,34.59,5335,0,Dos Palos,1,1,Fiber Optic,37.045728000000004,-120.63068200000001,0,74.9,0,0,Offer E,9388,0,0,0,0,7,0,0.0,242.13,0.0,490.55,0,1,93620
2448,0,1,0,0,14,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.85,1531.4,1,80,8,29.96,2292,1,Dunlap,1,0,Cable,36.789213000000004,-119.14033799999999,0,109.044,0,0,None,506,0,4,0,0,14,1,123.0,419.44,0.0,1531.4,0,0,93621
2449,1,0,1,1,11,1,0,DSL,0,0,1,0,Month-to-month,1,Bank transfer (automatic),59.65,683.25,0,25,47,21.14,2136,0,Firebaugh,1,1,Fiber Optic,36.785618,-120.625382,1,59.65,1,7,Offer D,9491,0,0,1,0,11,2,0.0,232.54,0.0,683.25,1,1,93622
2450,0,0,1,1,72,1,1,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),110.45,8058.85,0,62,14,46.63,4754,0,Fish Camp,1,0,Fiber Optic,37.483534999999996,-119.679414,1,110.45,1,9,None,77,1,0,1,1,72,0,0.0,3357.36,0.0,8058.85,0,1,93623
2451,1,0,1,1,28,1,1,Fiber optic,1,1,1,1,One year,0,Electronic check,106.1,2847.4,1,58,26,9.62,3770,1,Five Points,0,1,Fiber Optic,36.397745,-120.11991100000002,1,110.344,0,1,Offer C,1852,0,1,1,1,28,2,740.0,269.36,0.0,2847.4,0,0,93624
2452,1,1,0,0,15,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.2,1133.9,1,74,10,23.53,4553,1,Fowler,0,1,Fiber Optic,36.625792,-119.67248300000001,0,77.168,0,0,None,5635,0,2,0,0,15,4,0.0,352.9500000000001,43.31,1133.9,0,1,93625
2453,0,1,0,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.45,294.45,0,65,7,4.29,4093,0,Friant,0,0,DSL,37.027663000000004,-119.69056,0,74.45,0,0,None,1125,0,0,0,0,4,0,21.0,17.16,0.0,294.45,0,0,93626
2454,0,0,0,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,24.55,1719.15,0,30,0,2.66,4555,0,Helm,0,0,NA,36.520537,-120.118055,0,24.55,0,0,None,152,0,0,0,0,71,1,0.0,188.86,0.0,1719.15,0,0,93627
2455,0,0,0,0,5,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.35,461.7,1,30,76,10.11,4584,1,Hume,0,0,Fiber Optic,36.807595,-118.901544,0,92.924,0,0,Offer E,93,1,1,0,1,5,2,351.0,50.55,0.0,461.7,0,0,93628
2456,1,0,1,1,47,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.55,1160.45,0,28,0,15.68,3629,0,Kerman,0,1,NA,36.727418,-120.123526,1,24.55,2,3,Offer B,14062,0,0,1,0,47,0,0.0,736.96,0.0,1160.45,1,0,93630
2457,1,1,1,0,57,1,0,Fiber optic,0,1,1,0,One year,1,Electronic check,90.65,5199.8,0,66,4,46.62,5636,0,Kingsburg,1,1,Cable,36.478239,-119.52136999999999,1,90.65,0,10,None,14088,0,0,1,0,57,0,208.0,2657.34,0.0,5199.8,0,0,93631
2458,1,1,1,0,50,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),105.05,5163.3,0,77,8,40.9,5324,0,Lakeshore,1,1,Fiber Optic,37.290606,-119.216328,1,105.05,0,1,None,52,0,0,1,1,50,1,0.0,2045.0,0.0,5163.3,0,1,93634
2459,1,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.45,162.3,0,23,0,35.21,5624,0,Los Banos,0,1,NA,36.995162,-120.955099,0,20.45,0,0,Offer E,29124,0,0,0,0,8,1,0.0,281.68,0.0,162.3,1,0,93635
2460,0,0,1,1,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.55,883.35,0,20,0,13.26,5461,0,Madera,0,0,NA,36.902954,-120.194274,1,19.55,2,3,Offer B,28434,0,1,1,0,48,2,0.0,636.48,0.0,883.35,1,0,93637
2461,0,0,0,0,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.7,1341.5,0,30,0,10.0,6072,0,Madera,0,0,NA,37.004068,-119.930027,0,19.7,0,0,None,49247,0,0,0,0,70,1,0.0,700.0,0.0,1341.5,0,0,93638
2462,1,0,0,1,1,1,0,DSL,1,1,0,1,Month-to-month,1,Bank transfer (automatic),70.45,70.45,0,61,21,20.1,2706,0,Escondido,0,1,Cable,33.141265000000004,-116.967221,0,70.45,1,0,None,48690,1,0,0,1,1,1,0.0,20.1,0.0,70.45,0,1,92027
2463,1,0,1,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),85.65,659.45,0,62,16,39.59,2512,0,Miramonte,0,1,Fiber Optic,36.696759,-119.024051,1,85.65,0,1,Offer E,571,0,0,1,1,8,0,0.0,316.72,0.0,659.45,0,1,93641
2464,0,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,77.15,77.15,1,32,21,27.7,2756,1,North Fork,0,0,Cable,37.244307,-119.470256,0,80.236,0,0,None,3376,0,0,0,0,1,4,0.0,27.7,0.0,77.15,0,0,93643
2465,1,0,0,0,1,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Bank transfer (automatic),35.25,35.25,1,53,10,0.0,2548,1,Oakhurst,0,1,Cable,37.648647,-119.231447,0,36.66,0,0,None,8521,0,0,0,1,1,1,0.0,0.0,0.0,35.25,0,1,93644
2466,1,0,1,1,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.55,1205.05,0,37,0,15.65,4020,0,O Neals,0,1,NA,37.140104,-119.65709199999999,1,20.55,3,4,Offer B,173,0,1,1,0,60,2,0.0,939.0,0.0,1205.05,0,0,93645
2467,1,0,1,1,49,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,97.95,4917.9,0,61,18,16.02,4301,0,Orange Cove,0,1,DSL,36.633497999999996,-119.298895,1,97.95,1,7,Offer B,8449,1,0,1,1,49,1,88.52,784.98,0.0,4917.9,0,1,93646
2468,1,0,1,0,4,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,48.55,201,1,26,84,0.0,3955,1,Orosi,0,1,Fiber Optic,36.600184999999996,-119.175655,1,50.492,0,4,None,9780,0,2,1,1,4,4,169.0,0.0,0.0,201.0,1,0,93647
2469,0,0,0,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.0,599.3,0,30,0,32.43,4128,0,Parlier,0,0,NA,36.622237,-119.521126,0,20.0,0,0,Offer C,12587,0,0,0,0,29,0,0.0,940.47,0.0,599.3,0,0,93648
2470,0,0,1,0,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.25,1733.15,0,55,0,35.34,5887,0,Fresno,0,0,NA,36.841654999999996,-119.79711299999998,1,25.25,0,1,None,3258,0,0,1,0,67,0,0.0,2367.78,0.0,1733.15,0,0,93650
2471,0,0,1,0,53,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),98.4,5149.5,1,45,26,41.74,6481,1,Prather,0,0,Cable,37.007238,-119.505661,1,102.336,0,1,None,1314,0,0,1,1,53,5,133.89,2212.2200000000007,0.0,5149.5,0,1,93651
2472,1,0,1,0,67,1,1,DSL,1,1,0,0,Two year,0,Credit card (automatic),70.9,4677.1,0,38,15,28.06,4361,0,Raisin City,1,1,Cable,36.594542,-119.905245,1,70.9,0,8,None,265,1,0,1,0,67,1,70.16,1880.02,0.0,4677.1,0,1,93652
2473,0,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,119.3,0,40,0,6.48,5060,0,Raymond,0,0,NA,37.252057,-119.95783,1,19.85,1,1,Offer E,972,0,1,1,0,6,2,0.0,38.88,0.0,119.3,0,0,93653
2474,0,0,0,0,47,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.35,4849.1,0,51,10,14.54,3723,0,Reedley,1,0,Fiber Optic,36.636638,-119.421842,0,106.35,0,0,Offer B,25923,0,0,0,1,47,0,0.0,683.38,0.0,4849.1,0,1,93654
2475,0,0,0,0,53,1,0,Fiber optic,1,1,0,1,Two year,0,Mailed check,99.5,5424.25,0,46,13,43.57,4754,0,Riverdale,1,0,Cable,36.452211,-119.94575,0,99.5,0,0,Offer B,5729,1,0,0,1,53,0,0.0,2309.21,0.0,5424.25,0,1,93656
2476,1,0,1,0,69,1,0,DSL,1,1,1,1,Two year,1,Mailed check,84.7,5878.9,0,41,7,48.37,5345,0,Sanger,1,1,DSL,36.819628,-119.44041399999999,1,84.7,0,10,None,28991,1,0,1,1,69,0,412.0,3337.53,0.0,5878.9,0,0,93657
2477,1,0,0,0,3,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Mailed check,86.05,244.85,0,54,29,18.26,2500,0,San Joaquin,0,1,DSL,36.600193,-120.153393,0,86.05,0,0,Offer E,4318,0,0,0,1,3,1,71.0,54.78,0.0,244.85,0,0,93660
2478,1,0,0,0,4,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.55,220.75,0,38,29,30.07,2124,0,Selma,0,1,Fiber Optic,36.545322,-119.64228100000001,0,44.55,0,0,Offer E,26213,0,0,0,0,4,2,0.0,120.28,0.0,220.75,0,1,93662
2479,1,0,1,1,56,1,1,DSL,1,1,0,1,Two year,1,Credit card (automatic),75.85,4261.2,0,33,26,37.58,5314,0,Shaver Lake,0,1,Fiber Optic,37.223,-119.001021,1,75.85,1,6,Offer B,642,1,0,1,1,56,0,1108.0,2104.48,0.0,4261.2,0,0,93664
2480,1,1,1,0,59,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),93.85,5574.75,1,70,16,10.78,5390,1,South Dos Palos,0,1,DSL,36.959731,-120.65351899999999,1,97.604,0,0,None,343,0,1,0,0,59,3,892.0,636.02,8.13,5574.75,0,0,93665
2481,1,1,1,0,61,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.0,1501.75,0,68,0,19.14,6421,0,Sultana,0,1,NA,36.545353000000006,-119.33853500000001,1,25.0,0,5,None,306,0,0,1,0,61,1,0.0,1167.54,0.0,1501.75,0,0,93666
2482,0,0,1,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.0,89.75,0,38,12,15.5,5225,0,Tollhouse,0,0,Fiber Optic,36.993666,-119.34826699999999,1,45.0,0,8,Offer E,2633,0,0,1,0,2,1,0.0,31.0,0.0,89.75,0,1,93667
2483,1,1,1,1,46,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,100.7,4541.2,1,76,19,49.11,5712,1,Tranquillity,1,1,Fiber Optic,36.635661,-120.28864399999999,1,104.728,0,3,None,1130,0,2,1,0,46,3,86.28,2259.06,46.64,4541.2,0,1,93668
2484,1,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.5,255.5,0,57,0,46.06,2891,0,Wishon,0,1,NA,37.287758000000004,-119.548156,1,20.5,1,6,None,327,0,0,1,0,12,0,0.0,552.72,0.0,255.5,0,0,93669
2485,0,0,0,0,14,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,80.45,1072,1,44,25,1.19,4155,1,Traver,1,0,DSL,36.456091,-119.486225,0,83.66799999999999,0,0,None,646,0,1,0,0,14,1,0.0,16.66,0.0,1072.0,0,1,93673
2486,0,0,1,1,28,1,1,Fiber optic,0,0,0,1,One year,1,Electronic check,90.45,2509.25,0,44,19,26.28,5823,0,Squaw Valley,0,0,Fiber Optic,36.719141,-119.20267700000001,1,90.45,1,7,Offer C,3146,1,0,1,1,28,0,0.0,735.84,0.0,2509.25,0,1,93675
2487,1,0,0,0,24,1,0,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),60.45,1440.75,0,50,4,23.71,5095,0,Fresno,0,1,DSL,36.749403,-119.78757399999999,0,60.45,0,0,Offer C,13858,1,1,0,0,24,1,0.0,569.04,0.0,1440.75,0,1,93701
2488,1,0,0,0,31,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,55.25,1715.65,1,60,7,1.53,2933,1,Fresno,1,1,Cable,36.739385,-119.753649,0,57.46,0,0,Offer C,47999,1,0,0,0,31,5,120.0,47.43,0.0,1715.65,0,0,93702
2489,0,0,1,1,68,1,1,DSL,1,1,0,1,One year,1,Electronic check,78.45,5333.35,0,57,29,7.47,5071,0,Fresno,1,0,Fiber Optic,36.768774,-119.76263300000001,1,78.45,3,8,None,31180,1,0,1,1,68,1,154.67,507.96,0.0,5333.35,0,1,93703
2490,1,0,0,1,39,1,1,Fiber optic,0,0,1,1,Two year,0,Mailed check,100.55,3895.35,0,21,85,14.72,3124,0,Fresno,0,1,Fiber Optic,36.799648,-119.801247,0,100.55,1,0,Offer C,26580,1,0,0,1,39,1,0.0,574.08,0.0,3895.35,1,1,93704
2491,0,0,1,0,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.35,869.9,0,37,0,5.95,2127,0,Fresno,0,0,NA,36.787240000000004,-119.82781299999999,1,20.35,0,0,Offer B,35451,0,0,0,0,42,0,0.0,249.9,0.0,869.9,0,0,93705
2492,1,0,1,0,13,0,No phone service,DSL,1,0,1,1,Month-to-month,1,Electronic check,54.45,706.85,1,28,78,0.0,5212,1,Fresno,0,1,Fiber Optic,36.654614,-119.903674,1,56.62800000000001,0,1,None,35790,1,2,1,1,13,4,551.0,0.0,0.0,706.85,1,0,93706
2493,0,0,1,0,6,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,90.75,512.25,0,56,8,23.35,4297,0,Fresno,0,0,Fiber Optic,36.822715,-119.761826,1,90.75,0,1,None,29337,0,0,1,1,6,0,0.0,140.10000000000002,0.0,512.25,0,1,93710
2494,1,0,0,0,35,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),75.35,2636.05,1,53,23,25.04,2785,1,San Dimas,0,1,DSL,34.102119,-117.815532,0,78.36399999999998,0,0,Offer C,33878,0,0,0,0,35,2,606.0,876.4,0.0,2636.05,0,0,91773
2495,0,0,1,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.25,814.75,0,47,0,10.54,4411,0,Fresno,0,0,NA,36.878709,-119.7645,1,20.25,0,1,Offer C,45087,0,0,1,0,38,0,0.0,400.52,0.0,814.75,0,0,93720
2496,1,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.05,388.6,0,64,0,26.26,2782,0,Fresno,0,1,NA,36.732694,-119.783786,0,20.05,0,0,None,6848,0,0,0,0,18,2,0.0,472.68,0.0,388.6,0,0,93721
2497,0,0,1,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.6,93.45,0,34,0,29.14,4580,0,Fresno,0,0,NA,36.78979,-119.92989399999999,1,19.6,0,1,None,60889,0,0,1,0,4,0,0.0,116.56,0.0,93.45,0,0,93722
2498,1,0,1,0,27,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,53.8,1389.85,0,32,15,41.48,2563,0,Fresno,0,1,DSL,36.623632,-119.741322,1,53.8,0,1,Offer C,21010,1,0,1,0,27,0,0.0,1119.9599999999996,0.0,1389.85,0,1,93725
2499,1,0,0,1,41,1,0,DSL,1,1,1,0,One year,0,Mailed check,70.2,2894.55,0,44,11,13.76,5365,0,Fresno,1,1,DSL,36.793601,-119.761131,0,70.2,1,0,None,39148,0,0,0,0,41,0,0.0,564.16,0.0,2894.55,0,1,93726
2500,1,0,1,1,50,1,0,DSL,1,0,1,1,One year,0,Electronic check,75.5,4025.6,0,29,47,31.83,5141,0,Fresno,0,1,Fiber Optic,36.751489,-119.68072,1,75.5,1,1,None,54701,1,0,1,1,50,0,0.0,1591.5,0.0,4025.6,1,1,93727
2501,1,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,20.35,1354.4,0,24,0,22.78,4949,0,Fresno,0,1,NA,36.757345,-119.818274,1,20.35,1,1,None,16346,0,0,1,0,72,2,0.0,1640.16,0.0,1354.4,1,0,93728
2502,0,0,0,0,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),26.05,1856.4,0,35,0,31.33,4467,0,Salinas,0,0,NA,36.64152,-121.622188,0,26.05,0,0,None,35739,0,0,0,0,70,0,0.0,2193.1,0.0,1856.4,0,0,93901
2503,1,0,1,1,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.6,926,0,37,0,34.94,2471,0,Salinas,0,1,NA,36.667794,-121.60130600000001,1,20.6,2,1,None,58548,0,0,1,0,44,0,0.0,1537.36,0.0,926.0,0,0,93905
2504,1,0,0,0,2,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,75.7,189.2,1,55,2,42.16,4676,1,Salinas,0,1,Fiber Optic,36.722898,-121.633648,0,78.72800000000002,0,0,None,53946,0,2,0,0,2,1,0.38,84.32,0.0,189.2,0,1,93906
2505,0,0,1,1,34,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.1,682.1,0,43,0,41.72,2272,0,Salinas,0,0,NA,36.77462,-121.66471399999999,1,20.1,1,1,Offer C,22292,0,0,1,0,34,0,0.0,1418.48,0.0,682.1,0,0,93907
2506,0,1,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.3,1778.7,0,65,0,8.68,4397,0,Salinas,0,0,NA,36.624338,-121.615669,1,24.3,0,5,Offer A,13027,0,0,1,0,72,0,0.0,624.96,0.0,1778.7,0,0,93908
2507,1,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Electronic check,24.5,1816.2,0,20,0,32.18,4058,0,Escondido,0,1,NA,33.141265000000004,-116.967221,1,24.5,0,9,None,48690,0,0,1,0,71,0,0.0,2284.78,0.0,1816.2,1,0,92027
2508,0,0,0,0,64,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),110.5,7069.25,0,42,24,5.68,5718,0,Carmel By The Sea,1,0,Fiber Optic,36.554618,-121.92223899999999,0,110.5,0,0,None,2966,1,1,0,1,64,1,1697.0,363.52,0.0,7069.25,0,0,93921
2509,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.25,1841.2,0,45,0,49.51,4551,0,Carmel,0,0,NA,36.460611,-121.852507,1,25.25,0,9,None,13121,0,0,1,0,72,0,0.0,3564.72,0.0,1841.2,0,0,93923
2510,1,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.25,74.25,1,28,46,21.8,4750,1,Carmel Valley,0,1,Cable,36.414611,-121.6386,0,77.22,0,0,None,6691,0,0,0,0,1,0,0.0,21.8,0.0,74.25,1,0,93924
2511,1,1,1,0,29,1,0,Fiber optic,1,0,0,1,One year,0,Bank transfer (automatic),90.1,2656.7,0,73,16,32.03,3553,0,Chualar,1,1,Cable,36.596271,-121.442274,1,90.1,0,10,None,1140,0,0,1,1,29,2,425.0,928.87,0.0,2656.7,0,0,93925
2512,0,0,1,0,23,1,0,DSL,1,0,0,1,One year,1,Bank transfer (automatic),68.75,1689.45,0,38,29,31.39,3519,0,Gonzales,1,0,Fiber Optic,36.52588,-121.39671899999999,1,68.75,0,3,None,9023,1,0,1,1,23,1,0.0,721.97,0.0,1689.45,0,1,93926
2513,1,0,1,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.2,1054.75,0,19,0,40.76,4203,0,Greenfield,0,1,NA,36.248708,-121.38661699999999,1,19.2,3,10,None,14204,0,0,1,0,52,0,0.0,2119.52,0.0,1054.75,1,0,93927
2514,0,1,0,0,25,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.7,2187.55,1,72,7,36.36,4078,1,Jolon,0,0,Cable,35.930782,-121.189757,0,93.288,0,0,None,254,0,0,0,0,25,1,0.0,909.0,23.33,2187.55,0,1,93928
2515,0,0,0,0,64,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),115.1,7334.05,0,51,4,44.31,5213,0,King City,1,0,Cable,36.220760999999996,-120.980777,0,115.1,0,0,None,14477,1,0,0,1,64,0,29.34,2835.84,0.0,7334.05,0,1,93930
2516,0,1,0,0,16,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.4,1581.2,1,66,15,32.11,2688,1,Lockwood,0,0,Fiber Optic,35.989792,-121.05593300000001,0,100.256,0,0,None,538,0,0,0,0,16,2,237.0,513.76,47.2,1581.2,0,0,93932
2517,1,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.5,69.5,1,75,16,41.2,3273,1,Marina,0,1,Fiber Optic,36.689582,-121.758398,0,72.28,0,0,None,21759,0,0,0,0,1,2,0.0,41.2,0.0,69.5,0,1,93933
2518,1,0,0,0,24,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),99.65,2404.85,0,39,6,25.68,5207,0,Monterey,0,1,Cable,36.362741,-121.869685,0,99.65,0,0,Offer C,32857,0,0,0,1,24,1,144.0,616.3199999999998,0.0,2404.85,0,0,93940
2519,1,0,1,0,2,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,91.45,171.45,0,39,20,49.41,4889,0,Pacific Grove,1,1,Fiber Optic,36.618337,-121.92641699999999,1,91.45,0,0,None,15449,0,1,0,0,2,4,0.0,98.82,0.0,171.45,0,1,93950
2520,0,0,1,1,34,1,0,DSL,1,1,1,1,Two year,0,Mailed check,84.75,2839.45,0,41,16,9.09,2020,0,Pebble Beach,1,0,Fiber Optic,36.587497,-121.94481499999999,1,84.75,2,9,Offer C,4602,1,0,1,1,34,0,0.0,309.06,0.0,2839.45,0,1,93953
2521,1,1,1,0,36,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),85.25,3132.75,1,65,6,24.54,3041,1,San Lucas,0,1,Fiber Optic,36.125529,-120.864443,1,88.66,0,1,None,521,0,1,1,1,36,2,188.0,883.4399999999998,0.0,3132.75,0,0,93954
2522,1,0,1,1,53,1,1,DSL,0,0,1,1,One year,1,Mailed check,78.75,3942.45,0,43,56,31.86,5052,0,Seaside,1,1,Fiber Optic,36.625114,-121.82356499999999,1,78.75,3,7,None,38244,1,0,1,1,53,1,0.0,1688.58,0.0,3942.45,0,1,93955
2523,0,0,1,1,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.25,873.4,0,64,0,37.35,2070,0,Soledad,0,0,NA,36.414215999999996,-121.360597,1,20.25,1,8,None,13003,0,0,1,0,47,1,0.0,1755.45,0.0,873.4,0,0,93960
2524,1,0,0,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.9,1529.65,0,22,0,31.93,5730,0,Spreckels,0,1,NA,36.624641,-121.647195,0,19.9,1,0,None,407,0,0,0,0,72,1,0.0,2298.96,0.0,1529.65,1,0,93962
2525,1,0,1,1,72,1,1,Fiber optic,1,1,0,1,Two year,1,Credit card (automatic),97.75,6991.6,0,25,59,20.79,4054,0,Belmont,0,1,Fiber Optic,37.509366,-122.306132,1,97.75,3,1,None,25566,1,0,1,1,72,1,4125.0,1496.88,0.0,6991.6,1,0,94002
2526,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.4,19.4,1,52,0,3.14,4152,1,Brisbane,0,1,NA,37.684694,-122.40711999999999,0,19.4,0,0,None,3635,0,1,0,0,1,3,0.0,3.14,0.0,19.4,0,0,94005
2527,0,0,0,0,9,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,83.3,803.3,1,46,19,29.7,3520,1,Burlingame,0,0,DSL,37.57028,-122.365778,0,86.632,0,0,None,40346,0,0,0,1,9,3,153.0,267.3,0.0,803.3,0,0,94010
2528,0,0,0,0,8,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),80.1,679.3,1,34,8,36.39,5071,1,Daly City,0,0,Cable,37.691561,-122.445202,0,83.304,0,0,None,47453,0,3,0,0,8,1,0.0,291.12,0.0,679.3,0,1,94014
2529,1,1,0,0,45,1,0,DSL,1,0,0,1,One year,0,Credit card (automatic),62.7,2791.5,1,79,19,10.67,2654,1,Daly City,1,1,DSL,37.680844,-122.48131000000001,0,65.208,0,0,None,63337,0,0,0,0,45,6,0.0,480.15,0.0,2791.5,0,1,94015
2530,0,0,0,0,7,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.4,715,0,45,25,39.02,5041,0,Half Moon Bay,1,0,DSL,37.45567,-122.407992,0,100.4,0,0,None,17929,1,0,0,1,7,1,179.0,273.14000000000004,0.0,715.0,0,0,94019
2531,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.45,1681.6,0,59,0,33.0,4742,0,La Honda,0,0,NA,37.285677,-122.22416499999999,1,24.45,0,10,None,1622,0,0,1,0,71,3,0.0,2343.0,0.0,1681.6,0,0,94020
2532,0,1,0,0,41,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),101.1,4016.2,0,69,9,14.61,2227,0,Loma Mar,1,0,Cable,37.266388,-122.26308,0,101.1,0,0,None,148,1,0,0,1,41,0,0.0,599.01,0.0,4016.2,0,1,94021
2533,1,0,1,1,67,0,No phone service,DSL,1,0,1,1,Two year,0,Credit card (automatic),50.9,3281.65,0,39,17,0.0,5281,0,Los Altos,0,1,DSL,37.349546000000004,-122.13435600000001,1,50.9,2,2,Offer A,18486,0,0,1,1,67,0,558.0,0.0,0.0,3281.65,0,0,94022
2534,1,0,1,0,69,1,1,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),107.2,7317.1,0,51,24,33.37,5935,0,Los Altos,1,1,Fiber Optic,37.352911,-122.093002,1,107.2,0,8,Offer A,21496,1,0,1,1,69,1,0.0,2302.53,0.0,7317.1,0,1,94024
2535,0,1,1,0,70,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),92.2,6474.45,0,67,21,18.67,5264,0,Menlo Park,1,0,Cable,37.449551,-122.18376200000002,1,92.2,0,1,Offer A,39062,1,1,1,1,70,2,0.0,1306.9,0.0,6474.45,0,1,94025
2536,1,0,0,0,25,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),25.3,676.35,1,62,0,5.57,3779,1,Atherton,0,1,NA,37.454924,-122.20316799999999,0,25.3,0,0,Offer C,6876,0,0,0,0,25,6,0.0,139.25,0.0,676.35,0,0,94027
2537,1,0,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),113.4,8164.1,0,33,25,2.56,6347,0,Portola Valley,1,1,DSL,37.369709,-122.21584399999999,0,113.4,0,0,Offer A,6601,1,0,0,1,72,0,204.1,184.32,0.0,8164.1,0,1,94028
2538,1,0,1,1,34,0,No phone service,DSL,0,0,1,0,Two year,1,Electronic check,40.55,1325.85,0,31,29,0.0,3897,0,Millbrae,0,1,Fiber Optic,37.601248,-122.403099,1,40.55,1,10,None,20350,1,0,1,0,34,0,0.0,0.0,0.0,1325.85,0,1,94030
2539,0,0,1,1,65,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),26.0,1654.85,0,48,0,2.95,5352,0,Montara,0,0,NA,37.540582,-122.50959399999999,1,26.0,1,7,None,2346,0,0,1,0,65,0,0.0,191.75,0.0,1654.85,0,0,94037
2540,0,0,0,0,70,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),111.95,7795.95,0,60,26,44.57,4182,0,Moss Beach,1,0,Fiber Optic,37.515556,-122.502311,0,111.95,0,0,Offer A,3064,1,0,0,1,70,0,0.0,3119.9,0.0,7795.95,0,1,94038
2541,0,0,1,1,72,0,No phone service,DSL,1,0,1,1,Two year,1,Credit card (automatic),53.8,3952.45,0,61,14,0.0,4954,0,Mountain View,1,0,Fiber Optic,37.380662,-122.086022,1,53.8,1,10,Offer A,32143,0,0,1,1,72,1,553.0,0.0,0.0,3952.45,0,0,94040
2542,1,0,0,1,35,1,0,DSL,0,0,1,1,One year,1,Mailed check,72.1,2495.15,0,23,73,10.11,5510,0,Mountain View,0,1,Cable,37.388349,-122.075299,0,72.1,2,0,None,13483,1,0,0,1,35,2,182.15,353.85,0.0,2495.15,1,1,94041
2543,1,0,0,0,13,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Mailed check,98.15,1230.25,1,46,16,3.36,5525,1,Mountain View,0,1,DSL,37.419725,-122.062947,0,102.076,0,0,None,27822,0,1,0,1,13,3,197.0,43.68,0.0,1230.25,0,0,94043
2544,0,0,1,0,12,1,1,DSL,1,0,1,1,One year,0,Electronic check,78.85,876.75,0,46,17,25.09,2495,0,Pacifica,1,0,DSL,37.573633,-122.45516699999999,1,78.85,0,3,None,38885,0,1,1,1,12,2,0.0,301.08,0.0,876.75,0,1,94044
2545,0,0,1,1,62,1,0,DSL,1,0,1,0,One year,1,Bank transfer (automatic),70.75,4263.45,0,58,20,42.05,4133,0,Pescadero,1,0,Fiber Optic,37.22565,-122.297533,1,70.75,2,5,None,2055,1,0,1,0,62,2,853.0,2607.1,0.0,4263.45,0,0,94060
2546,0,0,0,0,25,1,0,DSL,1,0,1,1,Month-to-month,1,Credit card (automatic),76.15,1992.95,0,26,48,21.67,3955,0,Redwood City,0,0,Fiber Optic,37.461251000000004,-122.23541399999999,0,76.15,0,0,None,35737,1,0,0,1,25,2,957.0,541.75,0.0,1992.95,1,0,94061
2547,0,0,0,0,52,0,No phone service,DSL,1,1,0,0,Two year,0,Mailed check,39.1,1982.1,0,63,7,0.0,4247,0,Redwood City,0,0,Cable,37.410567,-122.297152,0,39.1,0,0,None,25569,1,0,0,0,52,2,13.87,0.0,0.0,1982.1,0,1,94062
2548,1,1,0,0,8,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),69.95,562.7,0,67,6,42.53,2939,0,Redwood City,0,1,DSL,37.499411,-122.19631799999999,0,69.95,0,0,None,32368,0,0,0,0,8,2,0.0,340.24,0.0,562.7,0,1,94063
2549,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,33.7,0,33,0,1.81,4978,0,Redwood City,0,1,NA,37.527497,-122.23094099999999,0,20.05,0,0,None,10658,0,0,0,0,2,0,0.0,3.62,0.0,33.7,0,0,94065
2550,0,0,1,1,56,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.05,1090.1,0,58,0,35.38,5172,0,San Bruno,0,0,NA,37.624435999999996,-122.43066100000001,1,20.05,3,10,None,39566,0,0,1,0,56,2,0.0,1981.28,0.0,1090.1,0,0,94066
2551,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.45,227.45,0,27,0,35.81,4862,0,San Carlos,0,0,NA,37.497915,-122.26736100000001,0,19.45,0,0,None,28098,0,0,0,0,12,1,0.0,429.72,0.0,227.45,1,0,94070
2552,0,0,1,0,47,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,26.9,1250.85,0,20,0,11.68,2382,0,San Gregorio,0,0,NA,37.331762,-122.341444,1,26.9,0,7,None,291,0,0,1,0,47,0,0.0,548.96,0.0,1250.85,1,0,94074
2553,1,1,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.2,37.2,0,80,0,7.03,4577,0,South San Francisco,0,1,NA,37.654436,-122.426468,0,19.2,0,0,None,60599,0,1,0,0,2,1,0.0,14.06,0.0,37.2,0,0,94080
2554,0,0,0,0,18,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.0,892.7,0,30,69,17.33,4952,0,Sunnyvale,1,0,Cable,37.378541,-122.02045600000001,0,50.0,0,0,None,64010,0,0,0,0,18,0,616.0,311.93999999999994,0.0,892.7,0,0,94086
2555,0,0,0,0,8,1,0,DSL,1,0,1,0,Month-to-month,1,Electronic check,60.0,487.75,0,43,24,46.78,5862,0,Sunnyvale,0,0,Cable,37.3511,-122.03731100000002,0,60.0,0,0,None,50070,0,1,0,0,8,1,117.0,374.24,0.0,487.75,0,0,94087
2556,1,0,1,0,45,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,84.55,3713.95,0,49,15,22.8,3289,0,Sunnyvale,1,1,Fiber Optic,37.421633,-122.00961299999999,1,84.55,0,8,None,16985,0,0,1,0,45,0,557.0,1026.0,0.0,3713.95,0,0,94089
2557,1,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.45,141.7,0,35,17,20.37,3666,0,San Francisco,0,1,Cable,37.7795,-122.419233,0,45.45,0,0,None,28998,0,0,0,0,3,1,2.41,61.11,0.0,141.7,0,1,94102
2558,0,0,0,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.05,678.2,0,22,0,40.64,4539,0,San Francisco,0,0,NA,37.773146999999994,-122.41128700000002,0,20.05,0,0,None,23036,0,0,0,0,38,0,0.0,1544.32,0.0,678.2,1,0,94103
2559,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,115.55,8425.3,0,46,21,47.82,5890,0,San Francisco,1,1,Cable,37.791222,-122.40224099999999,1,115.55,0,2,Offer A,384,1,1,1,1,72,2,0.0,3443.04,0.0,8425.3,0,1,94104
2560,1,0,0,0,46,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,93.7,4154.8,1,48,3,15.78,3378,1,San Francisco,0,1,Fiber Optic,37.789168,-122.395009,0,97.448,0,0,None,2066,0,1,0,1,46,3,125.0,725.88,0.0,4154.8,0,0,94105
2561,0,0,1,1,71,1,1,Fiber optic,1,1,1,0,Two year,1,Credit card (automatic),99.0,7061.65,0,43,17,15.73,4305,0,San Francisco,1,0,DSL,37.768881,-122.395521,1,99.0,2,4,Offer A,17372,0,0,1,0,71,2,0.0,1116.83,0.0,7061.65,0,1,94107
2562,1,0,1,1,66,0,No phone service,DSL,0,0,1,1,Two year,0,Bank transfer (automatic),50.55,3364.55,0,33,23,0.0,4652,0,San Francisco,0,1,Fiber Optic,37.791998,-122.408653,1,50.55,4,9,Offer A,13723,1,1,1,1,66,2,774.0,0.0,0.0,3364.55,0,0,94108
2563,1,1,0,0,25,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Mailed check,105.95,2655.25,1,73,24,46.34,4283,1,San Francisco,1,1,Cable,37.794487,-122.42227,0,110.18799999999999,0,0,Offer C,56330,0,2,0,0,25,2,637.0,1158.5,0.0,2655.25,0,0,94109
2564,1,0,0,0,18,1,1,DSL,0,0,1,1,One year,1,Credit card (automatic),82.0,1425.45,1,36,6,12.5,3306,1,San Francisco,1,1,Cable,37.750021000000004,-122.415201,0,85.28,0,0,None,74641,1,1,0,1,18,7,0.0,225.0,0.0,1425.45,0,1,94110
2565,0,0,1,1,13,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.0,332.5,0,44,0,35.19,4734,0,San Francisco,0,0,NA,37.801776000000004,-122.402293,1,25.0,3,5,None,3337,0,0,1,0,13,0,0.0,457.47,0.0,332.5,0,0,94111
2566,0,0,1,1,65,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),91.55,5963.95,0,52,26,10.11,4921,0,San Francisco,1,0,Fiber Optic,37.720498,-122.443119,1,91.55,3,1,None,73117,1,0,1,1,65,3,1551.0,657.15,0.0,5963.95,0,0,94112
2567,1,0,1,0,60,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,95.75,5742.9,1,59,18,35.22,4129,1,San Francisco,1,1,Cable,37.758084999999994,-122.43480100000001,1,99.58,0,1,None,30587,0,1,1,0,60,2,1034.0,2113.2,0.0,5742.9,0,0,94114
2568,1,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.35,278.85,0,19,0,46.47,2742,0,San Francisco,0,1,NA,37.786031,-122.437301,1,19.35,3,2,None,33122,0,1,1,0,15,2,0.0,697.05,0.0,278.85,1,0,94115
2569,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.85,1871.85,0,21,0,13.27,4067,0,San Francisco,0,0,NA,37.744409999999995,-122.486764,1,24.85,0,1,Offer A,42959,0,0,1,0,72,2,0.0,955.44,0.0,1871.85,1,0,94116
2570,1,0,1,0,30,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),94.05,2866.45,1,33,24,10.5,4095,1,San Francisco,0,1,Cable,37.770533,-122.445121,1,97.81200000000001,0,1,Offer C,38756,0,1,1,1,30,4,0.0,315.0,0.0,2866.45,0,1,94117
2571,0,0,1,1,42,1,0,Fiber optic,0,0,1,1,Two year,1,Electronic check,100.4,4303.65,0,42,26,12.6,3265,0,San Francisco,1,0,Fiber Optic,37.781304,-122.461522,1,100.4,3,1,None,38955,1,0,1,1,42,2,0.0,529.1999999999998,0.0,4303.65,0,1,94118
2572,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.0,1753,0,61,0,48.01,4066,0,San Francisco,0,0,NA,37.776718,-122.49578100000001,1,25.0,0,1,Offer A,42476,0,0,1,0,71,0,0.0,3408.71,0.0,1753.0,0,0,94121
2573,0,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,1,Mailed check,54.75,54.75,1,44,13,13.01,2614,1,San Francisco,0,0,Fiber Optic,37.760412,-122.48496599999999,0,56.94000000000001,0,0,None,55504,0,3,0,1,1,2,0.0,13.01,0.0,54.75,0,0,94122
2574,1,1,0,0,39,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.65,3759.05,1,79,25,41.93,4892,1,San Francisco,0,1,Fiber Optic,37.800253999999995,-122.436975,0,99.476,0,0,Offer C,22920,0,0,0,0,39,5,940.0,1635.27,0.0,3759.05,0,0,94123
2575,0,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.25,617.65,0,31,0,37.81,4988,0,San Francisco,0,0,NA,37.731505,-122.38453200000001,0,19.25,0,0,None,33177,0,0,0,0,35,0,0.0,1323.35,0.0,617.65,0,0,94124
2576,0,0,1,1,53,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),108.25,5935.1,0,38,29,43.39,5989,0,San Francisco,1,0,Cable,37.736534999999996,-122.45732,1,108.25,2,1,None,20643,1,2,1,1,53,2,1721.0,2299.67,0.0,5935.1,0,0,94127
2577,0,0,0,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.6,94.6,1,56,30,1.17,4033,1,San Francisco,0,0,Cable,37.797526,-122.46453100000001,0,98.384,0,0,None,2240,0,0,0,1,1,5,0.0,1.17,0.0,94.6,0,0,94129
2578,0,1,1,1,31,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.9,2911.3,1,70,23,47.95,4050,1,San Francisco,1,0,DSL,37.820894,-122.369725,1,102.856,0,1,Offer C,1458,1,0,1,0,31,4,0.0,1486.45,0.0,2911.3,0,1,94130
2579,1,0,0,0,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.15,982.95,0,41,0,33.68,4399,0,San Francisco,0,1,NA,37.746699,-122.44283300000001,0,20.15,0,0,None,27906,0,0,0,0,48,0,0.0,1616.64,0.0,982.95,0,0,94131
2580,0,1,0,1,30,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.3,2974.5,0,80,17,37.42,2440,0,San Francisco,0,0,DSL,37.722302,-122.491129,0,101.3,1,0,None,26297,1,0,0,1,30,0,0.0,1122.6,0.0,2974.5,0,1,94132
2581,1,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.0,198.7,0,56,0,4.42,2411,0,San Francisco,0,1,NA,37.802071000000005,-122.411004,0,20.0,0,0,None,26831,0,0,0,0,10,0,0.0,44.2,0.0,198.7,0,0,94133
2582,0,0,0,1,12,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.3,1275.65,0,62,18,16.96,5913,0,San Francisco,1,0,Fiber Optic,37.721052,-122.413573,0,105.3,2,0,None,40137,0,0,0,1,12,1,0.0,203.52,0.0,1275.65,0,1,94134
2583,0,1,0,0,57,1,0,DSL,1,0,1,0,Two year,0,Bank transfer (automatic),69.85,4003,0,67,30,11.23,4759,0,Palo Alto,1,0,Cable,37.444314,-122.149996,0,69.85,0,0,Offer B,16198,1,0,0,0,57,1,0.0,640.11,0.0,4003.0,0,1,94301
2584,0,0,1,0,58,1,0,DSL,1,1,1,0,Month-to-month,1,Credit card (automatic),65.25,3791.6,0,47,20,40.16,5912,0,Palo Alto,0,0,Cable,37.458090000000006,-122.115398,1,65.25,0,0,None,45499,0,0,0,0,58,1,0.0,2329.28,0.0,3791.6,0,1,94303
2585,0,0,0,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.8,813.3,0,49,0,41.99,5336,0,Palo Alto,0,0,NA,37.386978000000006,-122.177746,0,19.8,0,0,None,1723,0,0,0,0,37,0,0.0,1553.63,0.0,813.3,0,0,94304
2586,0,0,1,1,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.6,780.25,0,21,0,4.17,5584,0,Stanford,0,0,NA,37.424341999999996,-122.165641,1,19.6,2,1,None,13386,0,0,1,0,44,4,0.0,183.48,0.0,780.25,1,0,94305
2587,1,0,0,1,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.05,552.9,0,26,0,17.3,2400,0,Palo Alto,0,1,NA,37.416159,-122.13133700000002,0,20.05,3,0,None,24492,0,0,0,0,27,0,0.0,467.1,0.0,552.9,1,0,94306
2588,0,0,0,0,8,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,49.4,408.25,0,52,6,20.9,2907,0,San Mateo,0,0,DSL,37.590421,-122.306467,0,49.4,0,0,None,32488,1,0,0,0,8,0,2.45,167.2,0.0,408.25,0,1,94401
2589,1,1,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.05,231.8,1,71,31,30.25,2930,1,San Mateo,0,1,DSL,37.556634,-122.317723,0,79.092,0,0,None,23393,0,3,0,0,3,4,72.0,90.75,0.0,231.8,0,0,94402
2590,0,1,1,0,25,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Bank transfer (automatic),88.4,2191.15,0,72,4,19.44,4849,0,San Mateo,1,0,Fiber Optic,37.538309000000005,-122.305109,1,88.4,0,1,None,37926,0,0,1,1,25,2,0.0,486.00000000000006,0.0,2191.15,0,1,94403
2591,0,0,1,1,57,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.6,5611.7,0,37,28,32.37,6351,0,San Mateo,0,0,Fiber Optic,37.556094,-122.27243700000001,1,100.6,3,1,None,31882,0,0,1,1,57,0,0.0,1845.09,0.0,5611.7,0,1,94404
2592,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.45,246.25,0,38,0,18.12,4788,0,Alameda,0,0,NA,37.774633,-122.27443400000001,0,19.45,0,0,None,58555,0,0,0,0,12,2,0.0,217.44,0.0,246.25,0,0,94501
2593,0,0,1,1,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.3,1296.15,0,57,0,2.41,4574,0,Alameda,0,0,NA,37.724817,-122.22436299999998,1,20.3,2,1,None,13996,0,0,1,0,62,0,0.0,149.42000000000004,0.0,1296.15,0,0,94502
2594,0,0,1,0,65,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),107.65,7082.85,0,25,52,27.69,4193,0,Danville,1,0,DSL,37.791481,-121.903253,1,107.65,0,1,None,19777,1,0,1,1,65,1,0.0,1799.85,0.0,7082.85,1,1,94506
2595,0,0,1,0,71,1,1,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),80.45,5662.25,0,30,27,26.58,4518,0,Alamo,1,0,DSL,37.855717,-121.994813,1,80.45,0,1,Offer A,15187,1,0,1,1,71,0,0.0,1887.18,0.0,5662.25,0,1,94507
2596,0,0,1,1,21,1,0,DSL,0,1,1,0,One year,1,Credit card (automatic),58.85,1215.45,0,63,30,35.72,2845,0,Angwin,0,0,DSL,38.542448,-122.419923,1,58.85,3,1,None,3641,0,0,1,0,21,0,36.46,750.12,0.0,1215.45,0,1,94508
2597,1,0,1,0,71,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,109.6,7854.15,0,53,9,49.32,4564,0,Antioch,1,1,Fiber Optic,37.980057,-121.801599,1,109.6,0,9,Offer A,90891,0,0,1,1,71,0,70.69,3501.72,0.0,7854.15,0,1,94509
2598,0,0,0,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.15,525,0,56,10,30.06,4216,0,Benicia,1,0,DSL,38.113533000000004,-122.11926000000001,0,75.15,0,0,None,25578,0,0,0,0,7,0,0.0,210.42,0.0,525.0,0,1,94510
2599,0,0,0,0,72,1,0,DSL,1,1,0,1,Two year,1,Credit card (automatic),73.0,5265.2,0,23,69,23.02,5127,0,Bethel Island,1,0,Fiber Optic,38.050558,-121.646924,0,73.0,0,0,Offer A,2379,1,0,0,1,72,1,363.3,1657.44,0.0,5265.2,1,1,94511
2600,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.1,70.1,0,53,23,1.15,2475,0,Birds Landing,0,0,Fiber Optic,38.140719,-121.838298,0,70.1,0,0,None,138,0,0,0,0,1,0,0.0,1.15,0.0,70.1,0,1,94512
2601,0,0,1,1,72,1,1,Fiber optic,0,1,0,1,Two year,1,Bank transfer (automatic),98.65,7129.45,0,61,10,35.21,4616,0,Brentwood,1,0,Fiber Optic,37.908242,-121.682472,1,98.65,2,6,Offer A,26577,1,0,1,1,72,0,0.0,2535.12,0.0,7129.45,0,1,94513
2602,0,0,1,1,64,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,111.45,7266.95,0,48,53,39.37,5129,0,Byron,1,0,Fiber Optic,37.83323,-121.60146100000001,1,111.45,3,3,Offer B,10153,1,0,1,1,64,2,3851.0,2519.68,0.0,7266.95,0,0,94514
2603,0,0,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,114.9,8496.7,0,56,5,48.37,4589,0,Calistoga,1,0,DSL,38.629618,-122.593216,0,114.9,0,0,Offer A,7384,1,1,0,1,72,1,42.48,3482.64,0.0,8496.7,0,1,94515
2604,0,0,0,0,29,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),100.55,2878.75,0,33,12,10.67,4847,0,Clayton,1,0,Cable,37.881842,-121.84811100000002,0,100.55,0,0,None,14239,0,0,0,1,29,1,0.0,309.43,0.0,2878.75,0,1,94517
2605,0,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.4,261.3,0,23,0,6.56,4883,0,Concord,0,0,NA,37.950247999999995,-122.02245500000001,0,20.4,0,0,None,27394,0,0,0,0,13,1,0.0,85.28,0.0,261.3,1,0,94518
2606,0,0,0,0,31,1,1,Fiber optic,1,1,1,1,Month-to-month,0,Electronic check,104.35,3205.6,0,23,58,45.71,5320,0,Concord,0,0,DSL,37.990118,-122.012188,0,104.35,0,0,None,18650,0,0,0,1,31,1,1859.0,1417.01,0.0,3205.6,1,0,94519
2607,1,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.75,69.75,1,69,6,33.84,5057,1,Concord,0,1,Fiber Optic,38.013825,-122.039144,0,72.54,0,0,None,36186,0,3,0,0,1,3,0.0,33.84,0.0,69.75,0,1,94520
2608,1,0,1,1,7,0,No phone service,DSL,1,0,0,0,Month-to-month,1,Electronic check,34.5,279.25,1,61,33,0.0,3520,1,Concord,0,1,DSL,37.971421,-121.97150400000001,1,35.88,6,2,None,39888,1,5,1,0,7,4,0.0,0.0,0.0,279.25,0,1,94521
2609,1,0,1,0,61,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.55,6281.45,1,44,26,45.7,5011,1,Pleasant Hill,1,1,Cable,37.953379999999996,-122.07688600000002,1,109.772,0,1,None,32685,0,1,1,1,61,4,163.32,2787.7000000000007,0.0,6281.45,0,1,94523
2610,0,0,0,1,39,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),30.1,1131.3,1,56,26,0.0,3106,1,Crockett,1,0,Cable,38.049292,-122.22841499999998,0,31.304,2,0,None,3193,0,1,0,0,39,2,0.0,0.0,0.0,1131.3,0,1,94525
2611,1,0,1,0,10,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,738.2,1,36,25,31.72,2162,1,Danville,0,1,Fiber Optic,37.815459000000004,-121.977203,1,73.112,0,1,Offer D,32873,0,1,1,0,10,1,0.0,317.2,0.0,738.2,0,1,94526
2612,0,0,1,1,14,1,1,DSL,0,1,1,1,Month-to-month,0,Credit card (automatic),80.45,1137.05,0,43,21,9.77,5772,0,El Cerrito,0,0,DSL,37.924838,-122.28914499999999,1,80.45,3,8,Offer D,23141,1,0,1,1,14,1,239.0,136.78,0.0,1137.05,0,0,94530
2613,0,0,0,0,1,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,80.2,80.2,1,25,76,1.23,3056,1,Fairfield,0,0,Fiber Optic,38.287136,-122.02711000000001,0,83.40799999999999,0,0,Offer E,77683,0,0,0,0,1,4,0.0,1.23,0.0,80.2,1,0,94533
2614,0,0,1,1,67,1,1,Fiber optic,1,0,0,1,One year,1,Credit card (automatic),94.35,6341.45,1,41,12,30.94,4348,1,Travis Afb,0,0,Fiber Optic,38.265899,-121.93946100000001,1,98.124,0,1,Offer A,9978,1,1,1,1,67,3,76.1,2072.98,0.0,6341.45,0,1,94535
2615,0,0,0,0,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),91.35,6697.2,0,47,22,44.21,5378,0,Fremont,1,0,Cable,37.572272999999996,-121.964583,0,91.35,0,0,Offer A,66543,1,0,0,1,72,0,1473.0,3183.12,0.0,6697.2,0,0,94536
2616,1,0,1,1,6,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),44.6,260.8,1,61,23,49.2,4525,1,Fremont,0,1,Cable,37.505767999999996,-121.96247199999999,1,46.38399999999999,1,5,Offer E,56126,0,0,1,0,6,1,0.0,295.2000000000001,0.0,260.8,0,1,94538
2617,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.6,19.6,1,24,0,5.36,4205,1,Fremont,0,0,NA,37.516791,-121.89911699999999,0,19.6,0,0,Offer E,46917,0,0,0,0,1,4,0.0,5.36,0.0,19.6,1,0,94539
2618,1,0,1,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.9,505.45,0,47,0,18.87,4134,0,Hayward,0,1,NA,37.674002,-122.076796,1,19.9,1,0,None,60274,0,0,0,0,25,1,0.0,471.75,0.0,505.45,0,0,94541
2619,0,1,0,0,33,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,110.45,3655.45,1,70,28,17.24,3401,1,Hayward,1,0,Cable,37.656695,-122.04836100000001,0,114.868,0,0,Offer C,11147,1,0,0,1,33,0,1024.0,568.92,0.0,3655.45,0,0,94542
2620,1,0,0,0,18,1,0,DSL,1,0,1,0,Month-to-month,1,Electronic check,68.35,1299.8,0,22,48,48.68,5993,0,Hayward,1,1,Cable,37.639215,-122.037554,0,68.35,0,0,Offer D,72993,1,0,0,0,18,0,0.0,876.24,0.0,1299.8,1,1,94544
2621,1,0,1,0,71,1,0,DSL,0,1,1,1,Two year,1,Credit card (automatic),79.1,5564.85,0,21,27,28.02,5872,0,Hayward,1,1,Fiber Optic,37.62984,-122.120843,1,79.1,0,6,Offer A,27311,1,0,1,1,71,1,1503.0,1989.42,0.0,5564.85,1,0,94545
2622,1,1,1,1,28,1,1,DSL,0,0,0,0,One year,1,Electronic check,51.0,1381.8,0,73,21,4.71,5195,0,Castro Valley,0,1,Fiber Optic,37.708327000000004,-122.083473,1,51.0,2,1,None,41698,0,1,1,0,28,2,290.0,131.88,0.0,1381.8,0,0,94546
2623,0,0,0,1,2,1,1,Fiber optic,1,0,0,0,Month-to-month,0,Credit card (automatic),80.55,188.1,0,56,11,5.3,5346,0,Hercules,0,0,Fiber Optic,37.991259,-122.214945,0,80.55,1,0,None,22479,0,0,0,0,2,0,0.0,10.6,0.0,188.1,0,1,94547
2624,1,0,1,1,17,1,1,DSL,0,1,0,0,Month-to-month,1,Mailed check,66.7,1077.05,0,48,53,29.87,2814,0,Lafayette,1,1,Cable,37.907777,-122.12716100000002,1,66.7,3,1,Offer D,23996,1,0,1,0,17,0,0.0,507.79,0.0,1077.05,0,1,94549
2625,1,0,0,0,56,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,86.4,4922.4,0,32,13,37.15,4449,0,Livermore,0,1,DSL,37.571748,-121.65956200000001,0,86.4,0,0,Offer B,75929,0,0,0,0,56,0,0.0,2080.4,0.0,4922.4,0,1,94550
2626,0,0,1,0,60,0,No phone service,DSL,1,1,0,1,One year,0,Electronic check,50.05,2911.5,0,31,4,0.0,5493,0,Castro Valley,1,0,Fiber Optic,37.722727,-122.02157,1,50.05,0,7,Offer B,13212,0,0,1,1,60,0,116.0,0.0,0.0,2911.5,0,0,94552
2627,0,0,0,0,33,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.7,826.1,0,60,0,36.5,3378,0,Martinez,0,0,NA,38.014457,-122.11543200000001,0,25.7,0,0,None,46677,0,0,0,0,33,0,0.0,1204.5,0.0,826.1,0,0,94553
2628,0,0,0,0,1,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Mailed check,83.4,83.4,0,49,9,43.06,5960,0,Fremont,0,0,DSL,37.555473,-122.080312,0,83.4,0,0,None,33883,1,0,0,0,1,2,0.0,43.06,0.0,83.4,0,1,94555
2629,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),70.7,140.7,1,21,94,36.06,5317,1,Moraga,0,1,DSL,37.827946000000004,-122.10718500000002,0,73.528,0,0,None,16510,0,0,0,0,2,0,0.0,72.12,0.0,140.7,1,1,94556
2630,1,0,1,0,63,1,1,Fiber optic,1,0,0,0,Two year,1,Credit card (automatic),84.65,5377.8,0,52,7,12.96,4604,0,Napa,0,1,Cable,38.489789,-122.27011,1,84.65,0,8,Offer B,63947,1,0,1,0,63,1,376.0,816.48,0.0,5377.8,0,0,94558
2631,1,1,1,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.25,665.45,1,71,2,42.92,2487,1,Napa,1,1,DSL,38.232389000000005,-122.32494399999999,1,103.22,0,1,None,26894,0,0,1,1,7,1,13.0,300.44,0.0,665.45,0,0,94559
2632,0,0,0,0,55,1,0,DSL,0,1,0,1,Two year,1,Mailed check,64.75,3617.1,0,63,20,27.0,4634,0,Newark,1,0,Fiber Optic,37.504133,-122.032347,0,64.75,0,0,Offer B,42491,0,0,0,1,55,0,0.0,1485.0,0.0,3617.1,0,1,94560
2633,0,0,1,0,65,1,1,Fiber optic,1,1,1,0,One year,1,Bank transfer (automatic),100.15,6643.5,0,35,6,36.62,4915,0,Oakley,0,0,Fiber Optic,37.999406,-121.686241,1,100.15,0,8,Offer B,27607,1,0,1,0,65,3,0.0,2380.3,0.0,6643.5,0,1,94561
2634,1,0,1,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.8,84.8,1,21,56,37.83,2627,1,Orinda,0,1,DSL,37.873915999999994,-122.20522,1,88.19200000000001,0,1,Offer E,17964,1,2,1,0,1,3,0.0,37.83,0.0,84.8,1,0,94563
2635,1,0,0,0,63,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.25,1559.3,0,28,0,4.01,4530,0,Pinole,0,1,NA,37.996462,-122.29371599999999,0,25.25,0,0,Offer B,16717,0,1,0,0,63,2,0.0,252.63,0.0,1559.3,1,0,94564
2636,0,1,1,0,70,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),113.0,7987.6,0,74,14,46.2,4588,0,Pittsburg,1,0,Cable,38.006046999999995,-121.91683400000001,1,113.0,0,8,Offer A,78816,1,0,1,0,70,1,0.0,3234.0,0.0,7987.6,0,1,94565
2637,0,0,1,1,36,0,No phone service,DSL,1,0,0,0,Two year,0,Credit card (automatic),40.65,1547.35,0,19,71,0.0,2564,0,Pleasanton,1,0,Fiber Optic,37.633361,-121.86239499999999,1,40.65,3,5,None,36669,1,0,1,0,36,0,1099.0,0.0,0.0,1547.35,1,0,94566
2638,1,0,0,0,52,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),105.0,5426.85,1,21,56,49.29,4630,1,Pope Valley,1,1,Fiber Optic,38.672708,-122.40321899999999,0,109.2,0,0,None,494,1,2,0,1,52,4,3039.0,2563.08,0.0,5426.85,1,0,94567
2639,1,0,0,0,22,1,1,DSL,1,0,0,0,Month-to-month,1,Electronic check,54.45,1127.35,1,62,8,7.28,2445,1,Dublin,0,1,DSL,37.713926,-121.928425,0,56.62800000000001,0,0,Offer D,29636,0,0,0,0,22,5,0.0,160.16,0.0,1127.35,0,1,94568
2640,1,0,0,0,22,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),94.95,2142.8,0,37,18,48.07,4242,0,Port Costa,1,1,Cable,38.035707,-122.196821,0,94.95,0,0,Offer D,173,1,0,0,1,22,1,0.0,1057.54,0.0,2142.8,0,1,94569
2641,0,1,0,0,5,1,0,DSL,1,1,0,0,Month-to-month,0,Credit card (automatic),59.9,287.85,0,79,27,43.99,3662,0,Rio Vista,0,0,Fiber Optic,38.148862,-121.737696,0,59.9,0,0,None,5246,1,1,0,0,5,1,7.77,219.95,0.0,287.85,0,1,94571
2642,0,0,1,0,47,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.3,4045.65,1,40,25,44.26,3631,1,Rodeo,1,0,Cable,38.027218,-122.23463000000001,1,88.712,0,1,None,8506,0,0,1,1,47,4,1011.0,2080.22,0.0,4045.65,0,0,94572
2643,0,0,0,0,33,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,83.35,2757.85,1,51,33,20.29,5456,1,Saint Helena,0,0,DSL,38.581354,-122.296283,0,86.684,0,0,None,9423,0,0,0,1,33,2,910.0,669.5699999999998,0.0,2757.85,0,0,94574
2644,1,0,0,0,18,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),33.5,600,1,59,29,0.0,5474,1,Deer Park,1,1,DSL,38.554383,-122.474773,0,34.84,0,0,Offer D,223,0,2,0,0,18,3,174.0,0.0,0.0,600.0,0,0,94576
2645,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.8,19.8,0,50,0,11.96,3129,0,San Leandro,0,0,NA,37.717196,-122.15933799999999,0,19.8,0,0,None,41871,0,1,0,0,1,1,0.0,11.96,0.0,19.8,0,0,94577
2646,1,0,0,0,56,1,0,DSL,0,1,1,1,Two year,1,Credit card (automatic),81.8,4534.45,0,55,21,49.36,4399,0,San Leandro,1,1,DSL,37.704384000000005,-122.126703,0,81.8,0,0,Offer B,36568,1,1,0,1,56,1,95.22,2764.16,0.0,4534.45,0,1,94578
2647,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.0,40.9,0,40,0,43.27,2237,0,San Leandro,0,0,NA,37.687264,-122.15728,0,20.0,0,0,Offer E,19815,0,0,0,0,2,0,0.0,86.54,0.0,40.9,0,0,94579
2648,1,0,0,0,35,1,1,DSL,1,0,0,0,Month-to-month,1,Electronic check,59.6,2094.9,0,48,16,20.61,2187,0,San Lorenzo,1,1,Fiber Optic,37.676249,-122.132415,0,59.6,0,0,None,26240,0,0,0,0,35,0,0.0,721.35,0.0,2094.9,0,1,94580
2649,0,0,1,0,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.0,1584.8,0,44,0,6.81,5538,0,San Ramon,0,0,NA,37.766556,-121.97678400000001,1,25.0,0,5,Offer B,44078,0,0,1,0,64,1,0.0,435.84,0.0,1584.8,0,0,94583
2650,0,0,0,0,15,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),84.35,1302.65,0,44,4,6.22,3314,0,Suisun City,1,0,Cable,38.197907,-122.01725800000001,0,84.35,0,0,Offer D,39279,0,0,0,0,15,0,52.0,93.3,0.0,1302.65,0,0,94585
2651,1,0,0,0,24,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.35,2238.5,1,64,25,32.49,5546,1,Sunol,0,1,Cable,37.587494,-121.86285600000001,0,93.964,0,0,None,790,0,2,0,1,24,1,560.0,779.76,0.0,2238.5,0,0,94586
2652,1,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,0,Mailed check,55.55,55.55,0,23,48,33.32,2207,0,Union City,0,1,Fiber Optic,37.59485,-122.051521,0,55.55,0,0,Offer E,66472,0,0,0,1,1,3,0.0,33.32,0.0,55.55,1,1,94587
2653,0,0,1,1,70,1,0,DSL,1,0,1,1,Two year,0,Credit card (automatic),75.35,5437.75,0,35,53,39.53,6477,0,Pleasanton,0,0,Fiber Optic,37.685052,-121.91206100000001,1,75.35,3,9,Offer A,28568,1,1,1,1,70,3,2882.0,2767.1,0.0,5437.75,0,0,94588
2654,1,0,1,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.75,90.75,1,26,57,23.06,5460,1,Vallejo,0,1,Cable,38.161321,-122.271588,1,94.38,0,0,Offer E,42209,0,0,0,1,1,4,0.0,23.06,0.0,90.75,1,1,94589
2655,0,0,0,1,4,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Mailed check,89.6,365.65,1,64,22,36.76,4689,1,Vallejo,0,0,DSL,38.104704999999996,-122.24738700000002,0,93.184,0,0,Offer E,37218,0,1,0,0,4,3,80.0,147.04,0.0,365.65,0,0,94590
2656,0,0,0,0,39,1,0,DSL,0,0,0,1,One year,0,Electronic check,59.3,2209.15,0,62,17,6.77,5843,0,Vallejo,0,0,Cable,38.105733,-122.18633799999999,0,59.3,0,0,None,51665,1,0,0,1,39,2,376.0,264.03,0.0,2209.15,0,0,94591
2657,0,0,0,0,29,1,1,DSL,1,0,0,1,Month-to-month,1,Electronic check,66.1,1912.15,0,32,26,17.87,5590,0,Vallejo,0,0,DSL,38.093701,-122.27658899999999,0,66.1,0,0,None,159,0,0,0,1,29,2,497.0,518.23,0.0,1912.15,0,0,94592
2658,0,0,1,1,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,18.8,255.55,0,38,0,44.55,5751,0,Walnut Creek,0,0,NA,37.862128000000006,-122.075197,1,18.8,3,2,Offer D,18024,0,0,1,0,14,0,0.0,623.6999999999998,0.0,255.55,0,0,94595
2659,0,0,0,0,61,1,1,DSL,1,0,1,1,Two year,0,Credit card (automatic),86.45,5175.3,0,57,24,4.51,4471,0,Walnut Creek,1,0,Fiber Optic,37.900662,-122.05278200000001,0,86.45,0,0,Offer B,40917,1,1,0,1,61,2,0.0,275.11,0.0,5175.3,0,1,94596
2660,1,0,0,1,13,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),52.1,670.65,0,28,59,19.17,4929,0,Walnut Creek,0,1,Fiber Optic,37.916647999999995,-122.00848300000001,0,52.1,1,0,Offer D,26022,0,0,0,1,13,3,0.0,249.21000000000004,0.0,670.65,1,1,94598
2661,0,0,0,0,66,0,No phone service,DSL,1,1,0,0,Two year,1,Mailed check,47.4,3177.25,0,64,29,0.0,6435,0,Yountville,1,0,Fiber Optic,38.421458,-122.365048,0,47.4,0,0,Offer A,2873,1,0,0,0,66,0,921.0,0.0,0.0,3177.25,0,0,94599
2662,1,0,0,0,2,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,49.25,90.35,1,21,56,0.0,5775,1,Oakland,1,1,DSL,37.776523,-122.219268,0,51.22,0,0,Offer E,54876,0,0,0,1,2,1,51.0,0.0,0.0,90.35,1,0,94601
2663,0,0,1,0,59,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),109.15,6557.75,0,52,4,40.47,5186,0,Oakland,1,0,Fiber Optic,37.803883,-122.208417,1,109.15,0,7,Offer B,28900,0,0,1,1,59,1,26.23,2387.73,0.0,6557.75,0,1,94602
2664,1,0,1,1,62,1,1,Fiber optic,1,1,1,0,One year,1,Credit card (automatic),94.95,5791.85,0,19,59,15.76,4262,0,Oakland,0,1,DSL,37.739113,-122.175602,1,94.95,3,6,Offer B,31392,0,1,1,1,62,1,341.72,977.12,0.0,5791.85,1,1,94603
2665,1,1,1,0,33,1,0,Fiber optic,1,1,0,1,One year,1,Electronic check,93.55,3055.5,0,73,18,44.54,4414,0,Oakland,0,1,Fiber Optic,37.758019,-122.138678,1,93.55,0,10,None,42854,1,0,1,0,33,3,0.0,1469.82,0.0,3055.5,0,1,94605
2666,1,0,0,1,66,1,0,DSL,0,1,1,1,Two year,1,Credit card (automatic),79.5,5196.1,0,48,23,12.48,4285,0,Oakland,1,1,Cable,37.792489,-122.24431399999999,0,79.5,2,0,Offer A,41876,1,0,0,1,66,1,0.0,823.6800000000002,0.0,5196.1,0,1,94606
2667,0,0,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),115.05,8405,0,41,15,19.6,5905,0,Oakland,1,0,DSL,37.80707,-122.29740100000001,0,115.05,0,0,Offer A,21054,1,2,0,1,72,1,1261.0,1411.2,0.0,8405.0,0,0,94607
2668,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.75,19.75,1,43,0,11.91,2611,1,Emeryville,0,1,NA,37.83726,-122.287648,0,19.75,3,0,None,24589,0,0,0,0,1,3,0.0,11.91,0.0,19.75,0,0,94608
2669,0,0,0,0,19,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,95.15,1789.25,1,64,19,32.87,5830,1,Oakland,0,0,DSL,37.834340999999995,-122.26437,0,98.956,0,0,Offer D,21097,0,0,0,1,19,2,340.0,624.53,0.0,1789.25,0,0,94609
2670,0,0,1,1,51,1,1,Fiber optic,1,0,1,0,One year,1,Mailed check,95.15,5000.05,0,21,47,18.42,6492,0,Oakland,0,0,Fiber Optic,37.808731,-122.238708,1,95.15,1,2,Offer B,29964,1,0,1,1,51,1,2350.0,939.42,0.0,5000.05,1,0,94610
2671,1,0,0,0,63,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,105.4,6713.2,0,25,73,22.73,4551,0,Oakland,0,1,DSL,37.828416,-122.21600500000001,0,105.4,0,0,Offer B,36517,1,0,0,1,63,0,4901.0,1431.99,0.0,6713.2,1,0,94611
2672,1,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.1,562.6,0,31,0,33.4,3428,0,Oakland,0,1,NA,37.809014000000005,-122.26973899999999,0,20.1,0,0,None,11702,0,0,0,0,27,0,0.0,901.8,0.0,562.6,0,0,94612
2673,1,0,0,0,22,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),101.35,2317.1,1,44,21,10.33,4694,1,Oakland,0,1,Cable,37.84551,-122.23518100000001,0,105.404,0,0,Offer D,15438,0,1,0,1,22,3,0.0,227.26,0.0,2317.1,0,1,94618
2674,0,1,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,91.45,0,65,0,41.98,3460,0,Oakland,0,0,NA,37.787186,-122.14633,0,20.05,0,0,None,24518,0,0,0,0,4,0,0.0,167.92,0.0,91.45,0,0,94619
2675,1,0,1,1,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.7,828.85,0,59,0,32.02,5320,0,Oakland,0,1,NA,37.750553000000004,-122.197175,1,20.7,1,10,Offer B,30751,0,1,1,0,42,2,0.0,1344.84,0.0,828.85,0,0,94621
2676,0,0,0,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.35,617.35,0,28,0,21.19,4840,0,Berkeley,0,0,NA,37.866009000000005,-122.28622800000001,0,20.35,0,0,None,15638,0,0,0,0,29,0,0.0,614.51,0.0,617.35,1,0,94702
2677,0,0,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),70.05,266.9,1,46,21,12.58,3600,1,Berkeley,0,0,Cable,37.863843,-122.27568400000001,0,72.852,0,0,None,19763,0,3,0,0,4,1,56.0,50.32,0.0,266.9,0,0,94703
2678,1,0,0,0,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.7,625.05,0,62,0,24.57,3302,0,Berkeley,0,1,NA,37.871415999999996,-122.246597,0,19.7,0,0,None,21205,0,0,0,0,30,2,0.0,737.1,0.0,625.05,0,0,94704
2679,1,0,1,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.65,301.4,1,24,33,48.64,4013,1,Berkeley,0,1,Cable,37.858897999999996,-122.24051200000001,1,77.63600000000002,0,8,None,12448,0,2,1,0,4,5,0.0,194.56,0.0,301.4,1,1,94705
2680,1,0,1,1,71,1,0,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),85.45,6029.9,0,35,53,22.83,5394,0,Albany,1,1,Fiber Optic,37.890274,-122.29519199999999,1,85.45,3,9,Offer A,15882,1,1,1,1,71,1,0.0,1620.9299999999996,0.0,6029.9,0,1,94706
2681,1,0,1,0,46,0,No phone service,DSL,1,0,0,0,Two year,0,Credit card (automatic),40.4,1842.7,0,63,26,0.0,2519,0,Berkeley,1,1,Fiber Optic,37.897753,-122.27939099999999,1,40.4,0,6,Offer B,11889,1,0,1,0,46,0,0.0,0.0,0.0,1842.7,0,1,94707
2682,1,0,0,0,4,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.4,206.6,1,60,11,30.44,4399,1,Berkeley,0,1,Cable,37.897743,-122.263124,0,52.416000000000004,0,0,None,10737,0,1,0,0,4,3,23.0,121.76,0.0,206.6,0,0,94708
2683,0,0,0,0,7,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,79.65,604.7,1,61,20,40.32,4513,1,Berkeley,0,0,Fiber Optic,37.878554,-122.26608999999999,0,82.83600000000001,0,0,None,10147,0,0,0,0,7,3,121.0,282.24,0.0,604.7,0,0,94709
2684,1,0,0,0,69,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),105.2,7386.05,0,48,28,44.57,6247,0,Berkeley,0,1,Fiber Optic,37.872902,-122.30370800000001,0,105.2,0,0,Offer A,8157,1,0,0,1,69,0,0.0,3075.33,0.0,7386.05,0,1,94710
2685,0,0,1,0,72,1,1,Fiber optic,1,1,1,0,Two year,0,Bank transfer (automatic),100.65,7334.05,0,48,28,41.68,6380,0,Richmond,1,0,DSL,37.945288,-122.383941,1,100.65,0,10,Offer A,28450,0,0,1,0,72,0,0.0,3000.96,0.0,7334.05,0,1,94801
2686,1,1,0,0,19,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,79.85,1471.75,1,67,16,16.78,3715,1,El Sobrante,1,1,Cable,37.963995000000004,-122.288296,0,83.044,0,0,None,25399,0,1,0,0,19,2,235.0,318.82000000000005,0.0,1471.75,0,0,94803
2687,1,0,0,0,28,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,91.0,2626.15,0,26,59,45.24,2448,0,Richmond,1,1,Fiber Optic,37.921034000000006,-122.341798,0,91.0,0,0,None,39089,1,0,0,1,28,0,0.0,1266.72,0.0,2626.15,1,1,94804
2688,1,0,1,0,5,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,78.75,412.1,1,55,8,1.16,3401,1,Richmond,0,1,DSL,37.941456,-122.320968,1,81.9,0,1,None,13984,0,1,1,0,5,3,33.0,5.8,0.0,412.1,0,0,94805
2689,0,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),116.75,8277.05,0,79,16,14.75,5098,0,San Pablo,1,0,Fiber Optic,37.980269,-122.34263500000002,1,116.75,0,6,Offer A,55720,1,0,1,0,72,2,1324.0,1062.0,0.0,8277.05,0,0,94806
2690,1,1,1,1,8,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),80.45,583.45,1,67,2,26.99,3443,1,San Rafael,0,1,Cable,37.972662,-122.491452,1,83.66799999999999,0,2,None,40239,0,1,1,0,8,3,0.0,215.92,0.0,583.45,0,1,94901
2691,0,0,0,0,7,1,0,DSL,1,0,0,1,One year,1,Electronic check,59.1,369.25,0,32,17,6.83,4770,0,San Rafael,0,0,DSL,38.018065,-122.546024,0,59.1,0,0,None,28403,0,0,0,1,7,0,0.0,47.81,0.0,369.25,0,1,94903
2692,0,0,0,0,22,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.8,1049.05,0,64,11,31.53,4667,0,Greenbrae,0,0,Cable,37.946616999999996,-122.563571,0,49.8,0,0,Offer D,12010,0,0,0,0,22,1,0.0,693.6600000000002,0.0,1049.05,0,1,94904
2693,1,0,0,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.3,1414.8,0,57,0,45.75,4722,0,Belvedere Tiburon,0,1,NA,37.885628999999994,-122.46858,0,19.3,0,0,None,13065,0,0,0,0,72,1,0.0,3294.0,0.0,1414.8,0,0,94920
2694,1,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.65,169.75,0,58,0,26.17,4535,0,Bodega,0,1,NA,38.343282,-122.9755,1,19.65,3,6,Offer E,584,0,1,1,0,8,2,0.0,209.36,0.0,169.75,0,0,94922
2695,1,0,1,0,52,1,1,DSL,1,1,0,1,One year,1,Credit card (automatic),81.4,4354.45,0,64,24,41.34,4628,0,Bodega Bay,1,1,Fiber Optic,38.377165000000005,-123.037957,1,81.4,0,6,Offer B,1785,1,0,1,1,52,0,1045.0,2149.6800000000007,0.0,4354.45,0,0,94923
2696,0,0,0,0,68,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,38.9,2719.2,0,21,58,0.0,5278,0,Bolinas,1,0,Fiber Optic,37.943087,-122.72379,0,38.9,0,0,None,1573,1,0,0,0,68,1,0.0,0.0,0.0,2719.2,1,1,94924
2697,0,0,1,0,71,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),87.95,6365.35,0,46,30,9.06,4278,0,Corte Madera,1,0,Cable,37.924014,-122.51169399999999,1,87.95,0,7,None,9038,1,0,1,1,71,1,1910.0,643.26,0.0,6365.35,0,0,94925
2698,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,51.6,0,27,0,27.47,3300,0,Rohnert Park,0,1,NA,38.347190000000005,-122.697822,0,19.85,0,0,Offer E,42544,0,0,0,0,2,2,0.0,54.94,0.0,51.6,1,0,94928
2699,0,1,0,0,34,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,96.35,3190.25,0,79,13,14.23,5425,0,Dillon Beach,0,0,DSL,38.24458,-122.956268,0,96.35,0,0,None,330,1,0,0,0,34,0,415.0,483.82,0.0,3190.25,0,0,94929
2700,0,0,0,0,35,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,24.15,812.5,0,54,21,0.0,5097,0,Fairfax,0,0,DSL,37.971751,-122.611873,0,24.15,0,0,None,8486,0,0,0,0,35,0,0.0,0.0,0.0,812.5,0,1,94930
2701,0,0,1,1,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.1,1143.8,0,21,0,42.11,4376,0,Cotati,0,0,NA,38.326215000000005,-122.71874199999999,1,19.1,1,8,None,7936,0,0,1,0,61,0,0.0,2568.71,0.0,1143.8,1,0,94931
2702,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.0,44,0,62,17,13.4,2785,0,Forest Knolls,0,1,Fiber Optic,38.010092,-122.68944199999999,0,44.0,0,0,Offer E,1025,0,0,0,0,1,1,0.0,13.4,0.0,44.0,0,0,94933
2703,0,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.1,50.1,1,47,15,46.49,4778,1,Inverness,0,0,Cable,38.099323,-122.945723,0,52.104000000000006,0,0,None,1004,0,1,0,0,1,5,0.0,46.49,0.0,50.1,0,1,94937
2704,0,0,1,1,53,1,0,DSL,0,0,0,1,One year,0,Credit card (automatic),60.6,3297,0,29,59,31.99,4854,0,Lagunitas,1,0,Cable,38.021772,-122.691744,1,60.6,5,3,None,821,0,0,1,1,53,0,0.0,1695.47,0.0,3297.0,1,1,94938
2705,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.65,1887,0,37,0,12.58,5613,0,Larkspur,0,0,NA,37.937082000000004,-122.53236899999999,1,25.65,0,4,None,6773,0,0,1,0,72,1,0.0,905.76,0.0,1887.0,0,0,94939
2706,1,0,1,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,76.4,151.8,1,19,56,20.5,4340,1,Marshall,1,1,DSL,38.129308,-122.83481499999999,1,79.456,0,1,Offer E,406,0,3,1,0,2,1,85.0,41.0,0.0,151.8,1,0,94940
2707,1,0,0,0,3,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.7,293.65,1,28,80,32.76,3916,1,Mill Valley,1,1,Cable,37.901371000000005,-122.572024,0,102.648,0,0,Offer E,28727,1,0,0,1,3,0,235.0,98.28,0.0,293.65,1,0,94941
2708,0,1,0,0,13,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,100.8,1308.1,1,69,31,7.22,3269,1,Novato,0,0,Cable,38.135897,-122.56368300000001,0,104.83200000000001,0,0,Offer D,16429,0,1,0,0,13,6,406.0,93.86,0.0,1308.1,0,0,94945
2709,1,1,1,0,41,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,53.95,2215.4,0,65,9,0.0,3920,0,Nicasio,1,1,Fiber Optic,38.065359,-122.665566,1,53.95,0,8,Offer B,607,0,0,1,1,41,1,0.0,0.0,0.0,2215.4,0,1,94946
2710,0,0,1,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.4,482.8,0,44,0,35.86,3071,0,Novato,0,0,NA,38.112165999999995,-122.63438400000001,1,20.4,0,6,None,24741,0,0,1,0,24,0,0.0,860.64,0.0,482.8,0,0,94947
2711,0,0,1,1,28,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),90.1,2598.95,1,37,14,18.31,5958,1,Novato,0,0,Cable,38.067204,-122.524004,1,93.704,0,1,None,13361,0,1,1,1,28,8,364.0,512.68,0.0,2598.95,0,0,94949
2712,1,0,0,0,8,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,29.35,216.45,0,47,8,0.0,5369,0,Olema,0,1,DSL,38.052209000000005,-122.775567,0,29.35,0,0,Offer E,248,0,0,0,0,8,0,17.0,0.0,0.0,216.45,0,0,94950
2713,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.45,20.45,0,28,0,42.17,2184,0,Penngrove,0,1,NA,38.325599,-122.642352,0,20.45,0,0,Offer E,3777,0,0,0,0,1,0,0.0,42.17,0.0,20.45,1,0,94951
2714,0,0,0,0,54,1,1,Fiber optic,0,0,0,1,Two year,1,Bank transfer (automatic),95.1,5064.85,0,26,52,11.76,4825,0,Petaluma,1,0,Cable,38.237018,-122.77871999999999,0,95.1,0,0,None,31930,1,0,0,1,54,1,0.0,635.04,0.0,5064.85,1,1,94952
2715,1,0,0,0,41,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),25.25,996.45,0,23,0,41.21,3461,0,Petaluma,0,1,NA,38.235021,-122.557332,0,25.25,0,0,None,35419,0,0,0,0,41,2,0.0,1689.61,0.0,996.45,1,0,94954
2716,0,0,1,0,19,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.9,839.65,0,33,22,34.51,5842,0,Point Reyes Station,0,0,DSL,38.060264000000004,-122.830646,1,44.9,0,0,Offer D,1885,0,0,0,0,19,2,0.0,655.6899999999998,0.0,839.65,0,1,94956
2717,0,0,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),92.65,6733,0,35,19,30.0,6342,0,San Anselmo,1,0,DSL,37.99272,-122.575026,1,92.65,1,4,None,16849,1,0,1,1,72,2,0.0,2160.0,0.0,6733.0,0,1,94960
2718,1,0,0,0,62,0,No phone service,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),43.7,2618.3,0,21,51,0.0,5254,0,San Geronimo,1,1,Fiber Optic,38.004740000000005,-122.66371699999999,0,43.7,0,0,None,548,1,0,0,0,62,2,133.53,0.0,0.0,2618.3,1,1,94963
2719,0,1,1,1,56,1,0,DSL,1,0,1,1,Two year,1,Credit card (automatic),72.6,4084.35,0,78,19,5.93,6357,0,San Quentin,0,0,DSL,37.942551,-122.491642,1,72.6,1,8,Offer B,6448,1,0,1,0,56,1,0.0,332.08,0.0,4084.35,0,1,94964
2720,1,0,0,0,15,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,51.55,765.5,1,47,29,3.15,2087,1,Sausalito,0,1,Cable,37.848641,-122.51569199999999,0,53.611999999999995,0,0,Offer D,11213,0,0,0,0,15,6,222.0,47.25,0.0,765.5,0,0,94965
2721,1,1,0,0,10,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.25,793.55,1,75,20,7.51,3856,1,Stinson Beach,0,1,DSL,37.921137,-122.65756200000001,0,82.42,0,0,Offer D,781,0,1,0,0,10,2,0.0,75.1,0.0,793.55,0,1,94970
2722,1,0,1,1,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,18.95,613.95,0,39,0,35.39,4735,0,Tomales,0,1,NA,38.240769,-122.90104099999999,1,18.95,1,2,None,384,0,0,1,0,32,0,0.0,1132.48,0.0,613.95,0,0,94971
2723,1,0,0,0,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.5,402.85,0,31,0,32.89,5654,0,Valley Ford,0,1,NA,38.339996,-122.935056,0,20.5,0,0,Offer D,66,0,0,0,0,21,3,0.0,690.69,0.0,402.85,0,0,94972
2724,1,0,1,1,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.95,1244.8,0,28,0,47.96,4803,0,Woodacre,0,1,NA,38.005839,-122.638155,1,19.95,2,9,None,1449,0,0,1,0,62,1,0.0,2973.52,0.0,1244.8,1,0,94973
2725,0,0,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,24.5,46.4,0,34,5,0.0,5786,0,Alviso,0,0,DSL,37.449537,-121.994813,0,24.5,0,0,Offer E,2147,0,0,0,0,2,0,2.0,0.0,0.0,46.4,0,0,95002
2726,1,0,0,1,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.6,581.85,0,42,0,8.55,2924,0,Aptos,0,1,NA,37.013471,-121.877877,0,20.6,2,0,None,24227,0,0,0,0,27,0,0.0,230.85,0.0,581.85,0,0,95003
2727,1,0,0,0,5,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),94.85,462.8,1,44,21,40.15,5701,1,Aromas,0,1,Fiber Optic,36.878364000000005,-121.62978100000001,0,98.644,0,0,Offer E,3373,0,2,0,1,5,4,0.0,200.75,0.0,462.8,0,1,95004
2728,0,0,0,0,25,0,No phone service,DSL,1,1,1,1,One year,0,Electronic check,61.05,1540.2,0,31,9,0.0,3695,0,Ben Lomond,1,0,DSL,37.078873,-122.09038600000001,0,61.05,0,0,None,6407,0,0,0,1,25,2,139.0,0.0,0.0,1540.2,0,0,95005
2729,0,0,0,0,2,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.7,169.8,1,39,7,14.07,2187,1,Boulder Creek,0,0,Cable,37.171727000000004,-122.14296100000001,0,89.12799999999999,0,0,None,10520,0,0,0,1,2,4,12.0,28.14,0.0,169.8,0,0,95006
2730,1,0,0,0,49,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),106.65,5168.1,0,45,25,22.52,5154,0,Brookdale,0,1,Cable,37.106902000000005,-122.10000600000001,0,106.65,0,0,None,1007,1,1,0,1,49,1,0.0,1103.48,0.0,5168.1,0,1,95007
2731,0,0,0,0,63,1,1,Fiber optic,1,1,1,1,Month-to-month,0,Credit card (automatic),108.25,6780.1,0,46,16,5.17,5331,0,Campbell,1,0,Fiber Optic,37.279689000000005,-121.954567,0,108.25,0,0,None,44976,0,0,0,1,63,2,0.0,325.71,0.0,6780.1,0,1,95008
2732,0,0,0,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.4,94.5,0,51,0,30.79,4929,0,Capitola,0,0,NA,36.977025,-121.95286399999999,0,20.4,3,0,Offer E,9673,0,0,0,0,4,2,0.0,123.16,0.0,94.5,0,0,95010
2733,0,0,1,0,1,1,0,DSL,0,0,1,0,Month-to-month,1,Mailed check,55.3,55.3,0,27,82,36.69,2849,0,Castroville,0,0,Fiber Optic,36.784481,-121.759054,1,55.3,0,8,None,8582,0,0,1,0,1,0,0.0,36.69,0.0,55.3,1,0,95012
2734,1,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,208,0,46,0,28.62,4032,0,Cupertino,0,1,NA,37.306612,-122.080621,0,20.25,0,0,Offer D,54431,0,0,0,0,11,2,0.0,314.82,0.0,208.0,0,0,95014
2735,1,1,0,0,52,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),72.95,3829.75,0,75,11,42.19,4368,0,Davenport,0,1,Fiber Optic,37.114335,-122.23716200000001,0,72.95,0,0,Offer B,857,0,0,0,0,52,2,0.0,2193.88,0.0,3829.75,0,1,95017
2736,0,1,1,0,60,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,89.45,5294.6,0,70,19,24.68,4340,0,Felton,0,0,DSL,37.089110999999995,-122.06221299999999,1,89.45,0,6,Offer B,8728,0,0,1,0,60,0,0.0,1480.8,0.0,5294.6,0,1,95018
2737,1,0,0,0,64,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),104.65,6889.8,0,47,23,25.95,6443,0,Freedom,1,1,Fiber Optic,36.936228,-121.785559,0,104.65,0,0,None,4753,1,0,0,1,64,1,158.47,1660.8,0.0,6889.8,0,1,95019
2738,0,0,1,1,43,1,0,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),75.2,3254.35,0,30,59,29.98,3976,0,Gilroy,1,0,DSL,37.03889,-121.52895500000001,1,75.2,1,10,None,49968,0,0,1,1,43,1,1920.0,1289.14,0.0,3254.35,0,0,95020
2739,0,0,1,0,61,1,1,Fiber optic,0,0,1,1,One year,0,Bank transfer (automatic),101.15,6383.9,0,35,23,36.13,5177,0,Escondido,0,0,Fiber Optic,33.141265000000004,-116.967221,1,101.15,0,5,None,48690,1,0,1,1,61,1,1468.0,2203.9300000000007,0.0,6383.9,0,0,92027
2740,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.4,44.4,1,58,33,26.53,3204,1,Los Gatos,0,0,Cable,37.222842,-121.988727,0,46.176,0,0,Offer E,13290,0,0,0,0,1,2,0.0,26.53,0.0,44.4,0,0,95030
2741,1,1,0,0,5,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.5,477.7,1,67,7,45.72,2718,1,Los Gatos,0,1,DSL,37.233034,-121.947427,0,93.08,0,0,None,24443,0,0,0,0,5,2,3.34,228.6,0.0,477.7,0,1,95032
2742,1,0,0,0,66,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),68.75,4447.55,0,64,10,20.52,5454,0,Los Gatos,1,1,DSL,37.160194,-121.94561100000001,0,68.75,0,0,None,10172,1,1,0,0,66,1,0.0,1354.32,0.0,4447.55,0,1,95033
2743,1,0,1,0,67,1,0,Fiber optic,1,1,1,1,Two year,1,Electronic check,111.05,7321.05,0,51,29,46.89,6103,0,Milpitas,1,1,DSL,37.441931,-121.878502,1,111.05,0,8,None,62848,1,0,1,1,67,1,0.0,3141.63,0.0,7321.05,0,1,95035
2744,0,0,1,0,42,1,0,Fiber optic,0,0,1,1,Two year,1,Credit card (automatic),99.0,4135,0,54,17,1.31,4545,0,Morgan Hill,1,0,Fiber Optic,37.161544,-121.649371,1,99.0,0,9,None,41707,1,0,1,1,42,0,703.0,55.02,0.0,4135.0,0,0,95037
2745,1,1,1,0,1,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.05,86.05,1,66,25,38.78,4843,1,Moss Landing,0,1,Fiber Optic,36.863303,-121.781632,1,89.492,0,0,None,899,0,4,0,0,1,2,0.0,38.78,0.0,86.05,0,0,95039
2746,0,0,1,1,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,21.0,697.7,0,60,0,9.8,5225,0,Mount Hermon,0,0,NA,37.051165999999995,-122.05619399999999,1,21.0,3,3,Offer C,77,0,0,1,0,31,3,0.0,303.8,0.0,697.7,0,0,95041
2747,1,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.4,168.65,0,63,0,9.19,5873,0,Paicines,0,1,NA,36.525703,-120.952122,0,19.4,0,0,None,813,0,0,0,0,7,0,0.0,64.33,0.0,168.65,0,0,95043
2748,1,0,0,0,4,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,44.55,174.3,1,44,22,0.0,5605,1,San Juan Bautista,0,1,DSL,36.810567999999996,-121.503022,0,46.332,0,0,Offer E,3402,0,0,0,1,4,3,3.83,0.0,0.0,174.3,0,1,95045
2749,1,0,1,1,34,1,1,DSL,0,0,1,1,One year,0,Bank transfer (automatic),77.2,2753.8,0,23,52,5.39,3997,0,San Martin,1,1,Fiber Optic,37.084697,-121.606417,1,77.2,1,0,Offer C,5671,0,2,0,1,34,1,0.0,183.26,0.0,2753.8,1,1,95046
2750,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.45,69.25,0,33,0,2.78,2787,0,Santa Clara,0,1,NA,37.351214,-121.952417,0,19.45,0,0,None,36349,0,0,0,0,3,0,0.0,8.34,0.0,69.25,0,0,95050
2751,0,0,1,1,19,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,24.85,434.8,0,21,85,0.0,2958,0,Santa Clara,0,0,DSL,37.348129,-121.98468999999999,1,24.85,1,4,Offer D,52986,0,0,1,0,19,1,36.96,0.0,0.0,434.8,1,1,95051
2752,1,0,1,1,31,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),35.4,1077.5,1,41,25,0.0,2067,1,Santa Clara,0,1,Fiber Optic,37.393553999999995,-121.96511399999999,1,36.816,3,1,None,13031,1,0,1,0,31,2,269.0,0.0,0.0,1077.5,0,0,95054
2753,0,0,0,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Mailed check,95.65,95.65,1,45,10,32.33,3473,1,Santa Cruz,0,0,DSL,36.993451,-122.098858,0,99.476,0,0,Offer E,43192,0,0,0,1,1,1,0.0,32.33,0.0,95.65,0,0,95060
2754,1,0,0,0,3,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,41.35,107.25,0,32,25,0.0,5534,0,Santa Cruz,1,1,Fiber Optic,36.974575,-121.991149,0,41.35,0,0,None,36631,1,0,0,0,3,2,27.0,0.0,0.0,107.25,0,0,95062
2755,1,0,1,0,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.6,851.2,0,59,0,16.07,5092,0,Santa Cruz,0,1,NA,37.007882,-122.065975,1,19.6,0,3,None,4563,0,0,1,0,46,0,0.0,739.22,0.0,851.2,0,0,95064
2756,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.95,20.95,1,19,0,40.48,4285,1,Santa Cruz,0,0,NA,37.031403999999995,-121.98186499999998,0,20.95,0,0,None,8365,0,0,0,0,1,0,0.0,40.48,0.0,20.95,1,0,95065
2757,0,0,1,1,69,1,1,Fiber optic,1,0,0,0,One year,0,Bank transfer (automatic),84.45,5848.6,0,47,16,38.92,5629,0,Scotts Valley,1,0,Fiber Optic,37.070177,-122.010077,1,84.45,1,7,None,14574,0,0,1,0,69,2,0.0,2685.48,0.0,5848.6,0,1,95066
2758,1,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,109.8,0,31,0,7.83,5064,0,Saratoga,0,1,NA,37.257771999999996,-122.051824,0,20.25,0,0,None,30589,0,0,0,0,5,0,0.0,39.15,0.0,109.8,0,0,95070
2759,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.65,19.65,0,20,0,27.88,3625,0,Soquel,0,1,NA,37.023669,-121.94646100000001,0,19.65,0,0,None,9823,0,1,0,0,1,2,0.0,27.88,0.0,19.65,1,0,95073
2760,1,0,0,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.65,595.5,0,28,0,31.53,2194,0,Watsonville,0,1,NA,36.931653999999995,-121.75238300000001,0,20.65,0,0,Offer C,81141,0,0,0,0,26,0,0.0,819.78,0.0,595.5,1,0,95076
2761,0,1,0,0,10,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,34.7,329.8,1,67,4,0.0,3244,1,San Jose,0,0,Cable,37.34667,-121.91001899999999,0,36.088,0,0,Offer D,18197,0,2,0,0,10,1,13.0,0.0,0.0,329.8,0,0,95110
2762,1,0,0,0,25,1,0,Fiber optic,0,0,1,1,Two year,0,Bank transfer (automatic),99.3,2513.5,0,21,51,4.94,3847,0,San Jose,1,1,Cable,37.284265000000005,-121.827673,0,99.3,0,0,Offer C,57748,1,0,0,1,25,1,0.0,123.5,0.0,2513.5,1,1,95111
2763,1,0,1,1,64,1,0,Fiber optic,1,1,0,0,Month-to-month,0,Electronic check,81.05,5135.35,0,47,12,49.49,5168,0,San Jose,0,1,Fiber Optic,37.343827000000005,-121.883119,1,81.05,2,4,None,52334,0,0,1,0,64,0,0.0,3167.36,0.0,5135.35,0,1,95112
2764,1,0,1,1,30,1,1,DSL,1,1,0,0,Month-to-month,0,Electronic check,67.6,2000.2,0,31,19,48.04,4104,0,San Jose,1,1,Fiber Optic,37.333851,-121.891147,1,67.6,1,4,Offer C,561,1,0,1,0,30,0,0.0,1441.2,0.0,2000.2,0,1,95113
2765,1,0,0,0,13,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.15,931.75,0,53,10,39.17,4599,0,San Jose,0,1,Fiber Optic,37.350284,-121.852855,0,70.15,0,0,Offer D,51706,0,1,0,0,13,1,0.0,509.21,0.0,931.75,0,1,95116
2766,0,0,1,0,64,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,115.0,7396.15,0,37,29,46.44,5189,0,San Jose,1,0,DSL,37.311088,-121.961786,1,115.0,0,1,None,29914,1,0,1,1,64,1,0.0,2972.16,0.0,7396.15,0,1,95117
2767,0,0,0,1,46,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),84.8,3958.85,0,28,59,4.08,5756,0,San Jose,1,0,Fiber Optic,37.255479,-121.88983799999998,0,84.8,2,0,None,31926,1,0,0,0,46,1,2336.0,187.68,0.0,3958.85,1,0,95118
2768,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.7,260.9,0,57,0,36.65,3423,0,San Jose,0,0,NA,37.233226,-121.78809,0,19.7,0,0,Offer D,10155,0,0,0,0,12,1,0.0,439.8,0.0,260.9,0,0,95119
2769,0,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.75,297.3,1,54,0,39.84,2428,1,San Jose,0,0,NA,37.186141,-121.843554,0,19.75,0,0,Offer D,37090,0,0,0,0,15,1,0.0,597.6,0.0,297.3,0,0,95120
2770,1,0,1,1,17,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,92.55,1515.1,1,42,14,17.71,5775,1,San Jose,0,1,Fiber Optic,37.304681,-121.809955,1,96.25200000000001,0,1,Offer D,37127,0,0,1,1,17,2,212.0,301.07,0.0,1515.1,0,0,95121
2771,0,0,1,1,13,1,0,DSL,1,0,0,1,Month-to-month,1,Mailed check,63.15,816.8,0,40,25,39.2,5916,0,San Jose,1,0,Cable,37.32886,-121.83456699999999,1,63.15,3,3,None,59841,0,0,1,1,13,0,0.0,509.6,0.0,816.8,0,1,95122
2772,0,0,1,1,67,1,1,DSL,1,1,1,0,Two year,0,Credit card (automatic),74.0,4868.4,0,49,16,43.01,4188,0,San Jose,0,0,Cable,37.238758000000004,-121.828375,1,74.0,2,5,None,59632,1,1,1,0,67,3,0.0,2881.67,0.0,4868.4,0,1,95123
2773,1,0,1,0,24,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,29.1,688,0,25,51,0.0,4636,0,San Jose,1,1,Fiber Optic,37.257063,-121.92303700000001,1,29.1,0,4,Offer C,45257,0,0,1,0,24,1,351.0,0.0,0.0,688.0,1,0,95124
2774,1,0,0,0,6,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.05,288.35,0,37,13,23.01,3929,0,San Jose,0,1,Fiber Optic,37.294926000000004,-121.89476299999998,0,50.05,0,0,Offer E,46185,1,0,0,0,6,1,37.0,138.06,0.0,288.35,0,0,95125
2775,1,1,1,0,53,1,1,DSL,1,0,0,0,One year,1,Electronic check,60.05,3229.65,1,71,7,21.67,5271,1,San Jose,0,1,DSL,37.327069,-121.91681899999999,1,62.452,0,1,None,27023,1,0,1,0,53,3,0.0,1148.51,0.0,3229.65,0,1,95126
2776,1,1,1,0,16,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),74.3,1178.25,1,74,9,26.12,2076,1,San Jose,0,1,Cable,37.375156,-121.79586699999999,1,77.27199999999999,0,1,Offer D,60620,0,2,1,0,16,1,106.0,417.92,0.0,1178.25,0,0,95127
2777,1,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.0,185.4,0,27,0,39.39,2706,0,San Jose,0,1,NA,37.316146,-121.93628500000001,0,20.0,0,0,None,32804,0,0,0,0,10,0,0.0,393.9,0.0,185.4,1,0,95128
2778,0,0,0,0,13,1,0,Fiber optic,0,1,0,0,One year,1,Mailed check,74.65,966.25,0,39,15,42.62,4172,0,San Jose,0,0,Fiber Optic,37.305622,-122.000887,0,74.65,0,0,None,37570,0,0,0,0,13,2,0.0,554.06,0.0,966.25,0,1,95129
2779,1,0,0,0,9,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.35,758.6,1,28,64,49.14,2752,1,San Jose,0,1,Cable,37.277592,-121.98647700000001,0,88.764,0,0,Offer E,13481,0,0,0,0,9,0,0.0,442.26,0.0,758.6,1,1,95130
2780,0,0,0,0,25,1,0,DSL,1,1,1,0,One year,0,Mailed check,74.3,1863.8,1,48,23,1.37,5175,1,San Jose,1,0,Cable,37.387027,-121.897775,0,77.27199999999999,0,0,None,26389,1,2,0,0,25,3,0.0,34.25,0.0,1863.8,0,1,95131
2781,1,1,0,0,7,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Electronic check,44.4,265.8,0,75,26,0.0,3410,0,San Jose,0,1,DSL,37.424655,-121.74841,0,44.4,0,0,None,40568,1,0,0,0,7,0,69.0,0.0,0.0,265.8,0,0,95132
2782,1,0,1,1,38,1,1,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),85.4,3297,0,26,59,17.52,5292,0,San Jose,1,1,Fiber Optic,37.371862,-121.860349,1,85.4,2,6,Offer C,26032,1,0,1,1,38,1,194.52,665.76,0.0,3297.0,1,1,95133
2783,0,0,1,0,43,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,94.1,4107.3,0,33,11,49.48,4392,0,San Jose,0,0,Fiber Optic,37.42765,-121.945416,1,94.1,0,9,None,9657,0,1,1,1,43,1,452.0,2127.64,0.0,4107.3,0,0,95134
2784,0,0,0,1,4,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),98.1,396.3,1,34,20,5.63,2895,1,San Jose,1,0,Cable,37.28682,-121.723877,0,102.024,0,0,Offer E,15798,1,0,0,1,4,5,79.0,22.52,0.0,396.3,0,0,95135
2785,0,0,0,0,25,1,1,Fiber optic,0,1,1,1,Two year,0,Electronic check,108.9,2809.05,0,20,51,32.33,4398,0,San Jose,1,0,DSL,37.270938,-121.851046,0,108.9,0,0,Offer C,36944,1,1,0,1,25,1,0.0,808.25,0.0,2809.05,1,1,95136
2786,1,0,0,1,27,1,0,DSL,1,1,0,0,One year,0,Mailed check,56.2,1567.55,0,19,59,2.63,5978,0,San Jose,0,1,DSL,37.246064000000004,-121.749494,0,56.2,2,0,Offer C,14792,0,1,0,0,27,1,925.0,71.00999999999998,0.0,1567.55,1,0,95138
2787,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,26.1,1851.45,0,61,0,33.92,5475,0,San Jose,0,1,NA,37.218705,-121.762429,1,26.1,2,2,None,7023,0,0,1,0,72,1,0.0,2442.24,0.0,1851.45,0,0,95139
2788,1,0,0,1,71,1,1,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),85.45,6028.95,0,19,30,31.89,4777,0,Mount Hamilton,0,1,Cable,37.382909000000005,-121.634151,0,85.45,1,0,None,38,0,0,0,0,71,0,1809.0,2264.19,0.0,6028.95,1,0,95140
2789,0,0,0,0,24,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),88.95,2072.75,0,63,9,44.09,5557,0,San Jose,1,0,Cable,37.339533,-121.777179,0,88.95,0,0,Offer C,44103,0,1,0,0,24,1,0.0,1058.16,0.0,2072.75,0,1,95148
2790,0,0,0,0,50,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,109.65,5551.15,1,63,31,27.7,5855,1,Stockton,0,0,Fiber Optic,37.959706,-121.287669,0,114.03600000000002,0,0,None,7071,1,0,0,1,50,0,1721.0,1385.0,0.0,5551.15,0,0,95202
2791,1,0,0,0,57,1,0,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),74.35,4317.35,0,30,42,24.67,5548,0,Stockton,1,1,Fiber Optic,37.954089,-121.329761,0,74.35,0,0,None,16357,0,0,0,1,57,0,0.0,1406.19,0.0,4317.35,0,1,95203
2792,0,0,0,0,15,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,48.85,736.8,0,34,23,31.68,5584,0,Stockton,0,0,Fiber Optic,37.974498,-121.31956799999999,0,48.85,0,0,None,30476,0,0,0,0,15,0,169.0,475.2,0.0,736.8,0,0,95204
2793,1,0,0,0,4,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,80.1,336.15,0,27,82,44.16,2333,0,Stockton,0,1,Fiber Optic,37.965695000000004,-121.260051,0,80.1,0,0,Offer E,34138,0,0,0,0,4,3,276.0,176.64,0.0,336.15,1,0,95205
2794,0,0,0,0,28,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,56.05,1522.65,0,51,15,44.11,4468,0,Stockton,0,0,Fiber Optic,37.902421999999994,-121.44002900000001,0,56.05,0,0,Offer C,49657,0,0,0,0,28,1,0.0,1235.08,0.0,1522.65,0,1,95206
2795,0,1,0,0,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.55,622.9,1,70,30,17.56,3145,1,Stockton,0,0,DSL,38.002125,-121.324979,0,77.532,0,0,None,49965,0,1,0,0,9,2,187.0,158.04,33.25,622.9,0,0,95207
2796,0,0,1,0,55,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Bank transfer (automatic),89.8,4959.6,0,37,9,5.08,5875,0,Stockton,0,0,Cable,38.044523,-121.34804799999999,1,89.8,0,2,Offer B,30814,0,0,1,0,55,1,446.0,279.4,0.0,4959.6,0,0,95209
2797,1,0,0,0,3,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.95,329.95,1,32,33,11.94,5351,1,Stockton,1,1,DSL,38.033219,-121.29743300000001,0,104.988,0,0,Offer E,40611,0,3,0,1,3,7,109.0,35.82,0.0,329.95,0,0,95210
2798,1,0,0,0,10,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.9,1048.85,1,25,45,40.22,2832,1,Stockton,1,1,Fiber Optic,38.049457000000004,-121.21653,0,98.696,0,0,Offer D,6951,0,3,0,1,10,7,472.0,402.2,0.0,1048.85,1,0,95212
2799,1,0,0,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.1,1001.5,0,53,0,39.29,4391,0,Stockton,0,1,NA,37.946282000000004,-121.139499,0,19.1,2,0,Offer B,23789,0,0,0,0,55,1,0.0,2160.95,0.0,1001.5,0,0,95215
2800,0,0,1,1,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,442.6,0,58,0,42.46,2522,0,Stockton,0,0,NA,38.029728999999996,-121.387999,1,20.35,3,9,None,19109,0,0,1,0,20,0,0.0,849.2,0.0,442.6,0,0,95219
2801,0,0,1,1,62,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),106.05,6703.5,0,47,23,15.05,6361,0,Acampo,0,0,Fiber Optic,38.200231,-121.23503400000001,1,106.05,2,8,Offer B,6317,1,0,1,1,62,1,1542.0,933.1,0.0,6703.5,0,0,95220
2802,1,1,1,0,32,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,104.9,3351.55,1,76,24,43.51,3966,1,Angels Camp,1,1,Cable,38.071327000000004,-120.632221,1,109.096,0,1,Offer C,4264,1,0,1,0,32,4,804.0,1392.32,33.73,3351.55,0,0,95222
2803,0,0,0,0,43,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.65,779.25,0,44,0,6.71,3678,0,Arnold,0,0,NA,38.321529999999996,-120.23635800000001,0,19.65,0,0,Offer B,5159,0,0,0,0,43,0,0.0,288.53,0.0,779.25,0,0,95223
2804,1,0,1,0,9,0,No phone service,DSL,0,0,0,0,One year,0,Bank transfer (automatic),24.1,259.8,1,53,16,0.0,3195,1,Avery,0,1,Cable,38.208335999999996,-120.33993799999999,1,25.064000000000004,0,1,Offer E,115,0,1,1,0,9,2,42.0,0.0,0.0,259.8,0,0,95224
2805,0,0,1,0,60,1,0,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),59.85,3483.45,0,49,21,41.4,4029,0,Burson,0,0,Fiber Optic,38.183918,-120.898817,1,59.85,0,7,Offer B,27,1,0,1,0,60,0,732.0,2484.0,0.0,3483.45,0,0,95225
2806,1,0,1,0,58,1,1,DSL,1,1,1,1,Two year,1,Electronic check,86.1,4890.5,0,38,2,22.14,5666,0,Campo Seco,1,1,Fiber Optic,38.233878999999995,-120.86166599999999,1,86.1,0,3,Offer B,75,0,1,1,1,58,2,0.0,1284.12,0.0,4890.5,0,1,95226
2807,1,0,0,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.45,136.75,0,47,0,49.16,5084,0,Clements,0,1,NA,38.227284999999995,-121.02788999999999,0,19.45,2,0,None,722,0,0,0,0,7,0,0.0,344.12,0.0,136.75,0,0,95227
2808,1,0,1,1,2,1,0,Fiber optic,1,0,1,1,Month-to-month,0,Electronic check,97.1,184.15,0,40,24,39.35,5745,0,Copperopolis,0,1,DSL,37.943954,-120.67108,1,97.1,1,10,Offer E,2633,0,1,1,1,2,3,0.0,78.7,0.0,184.15,0,1,95228
2809,1,1,0,0,37,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,36.65,1315,0,75,29,0.0,2494,0,Farmington,1,1,DSL,37.956963,-120.863055,0,36.65,0,0,Offer C,596,0,0,0,0,37,0,381.0,0.0,0.0,1315.0,0,0,95230
2810,0,1,1,1,65,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),103.9,6767.1,0,76,27,1.58,5669,0,French Camp,1,0,DSL,37.873283,-121.29203400000002,1,103.9,3,8,Offer B,5094,1,0,1,0,65,0,1827.0,102.7,0.0,6767.1,0,0,95231
2811,0,0,1,1,39,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,757.95,0,40,0,15.91,3944,0,Glencoe,0,0,NA,38.358464,-120.57930400000001,1,19.75,3,6,Offer C,21,0,0,1,0,39,0,0.0,620.49,0.0,757.95,0,0,95232
2812,1,0,1,0,66,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,104.05,6890,1,23,94,20.07,5504,1,Hathaway Pines,0,1,Cable,38.184914,-120.364085,1,108.212,0,1,Offer A,335,1,0,1,1,66,4,6477.0,1324.62,0.0,6890.0,1,0,95233
2813,1,0,0,0,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.55,1657.4,0,20,0,5.84,6042,0,Linden,0,1,NA,38.047746000000004,-121.030499,0,24.55,0,0,None,3148,0,0,0,0,68,2,0.0,397.12,0.0,1657.4,1,0,95236
2814,0,0,1,1,62,0,No phone service,DSL,1,1,1,0,Two year,0,Bank transfer (automatic),48.7,3008.55,0,32,26,0.0,5453,0,Lockeford,0,0,Cable,38.166790999999996,-121.14206999999999,1,48.7,2,6,Offer B,3205,1,0,1,0,62,0,0.0,0.0,0.0,3008.55,0,1,95237
2815,1,0,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,88.35,262.05,1,33,11,49.4,5202,1,Lodi,1,1,Cable,38.123544,-121.15907800000001,0,91.884,0,0,Offer E,45755,1,0,0,0,3,2,0.0,148.2,0.0,262.05,0,1,95240
2816,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,109.55,8165.1,0,34,2,44.2,6452,0,Lodi,1,0,Fiber Optic,38.128087,-121.4078,1,109.55,0,9,None,22073,0,0,1,1,72,1,163.0,3182.4,0.0,8165.1,0,0,95242
2817,0,0,1,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.65,875.55,0,40,0,8.44,5062,0,Mokelumne Hill,0,0,NA,38.304194,-120.592431,1,20.65,0,9,Offer B,2718,0,1,1,0,41,1,0.0,346.04,0.0,875.55,0,0,95245
2818,1,0,1,1,29,1,0,Fiber optic,1,0,1,1,Month-to-month,0,Credit card (automatic),94.65,2649.15,1,43,16,40.49,5150,1,Mountain Ranch,0,1,Fiber Optic,38.264262,-120.515133,1,98.436,0,1,None,1692,0,1,1,1,29,1,424.0,1174.21,0.0,2649.15,0,0,95246
2819,0,0,0,0,4,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,55.2,220.65,0,64,17,7.49,4042,0,Murphys,0,0,Cable,38.147852,-120.440124,0,55.2,0,0,Offer E,4353,0,0,0,0,4,0,38.0,29.96,0.0,220.65,0,0,95247
2820,1,0,0,0,53,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),24.05,1301.9,0,34,0,39.37,4865,0,San Andreas,0,1,NA,38.196496999999994,-120.61688999999998,0,24.05,0,0,Offer B,3930,0,0,0,0,53,0,0.0,2086.61,0.0,1301.9,0,0,95249
2821,1,1,1,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.4,74.4,1,67,32,17.36,5429,1,Sheep Ranch,0,1,Cable,38.244806,-120.417301,1,77.376,0,1,None,88,0,0,1,0,1,0,0.0,17.36,0.0,74.4,0,0,95250
2822,0,0,1,1,41,1,1,DSL,1,1,0,1,Month-to-month,0,Credit card (automatic),79.9,3326.2,1,42,62,45.26,4734,1,Vallecito,1,0,Fiber Optic,38.055562,-120.456298,1,83.096,3,1,None,460,1,2,1,1,41,3,2062.0,1855.66,0.0,3326.2,0,0,95251
2823,1,0,1,0,39,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.45,790,0,39,0,36.39,2165,0,Valley Springs,0,1,NA,38.156971,-120.849231,1,20.45,0,10,Offer C,11266,0,0,1,0,39,0,0.0,1419.21,0.0,790.0,0,0,95252
2824,1,0,1,0,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.25,1237.65,0,57,0,17.38,4538,0,Wallace,0,1,NA,38.192608,-120.957842,1,19.25,0,9,Offer B,304,0,1,1,0,63,1,0.0,1094.9399999999996,0.0,1237.65,0,0,95254
2825,1,0,0,0,15,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,26.35,378.6,0,48,0,7.96,2723,0,West Point,0,1,NA,38.41935,-120.469545,0,26.35,0,0,None,2198,0,1,0,0,15,2,0.0,119.4,0.0,378.6,0,0,95255
2826,0,0,1,0,13,1,0,DSL,0,0,0,0,One year,0,Electronic check,43.8,592.65,0,34,2,29.49,4369,0,Wilseyville,0,0,Cable,38.392686,-120.415951,1,43.8,0,1,None,435,0,0,1,0,13,0,12.0,383.37,0.0,592.65,0,0,95257
2827,1,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,50.15,50.15,0,45,16,20.3,4014,0,Woodbridge,0,1,DSL,38.169605,-121.31096399999998,0,50.15,0,0,Offer E,4176,0,0,0,0,1,1,0.0,20.3,0.0,50.15,0,0,95258
2828,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.45,20.45,0,37,0,43.82,5925,0,Atwater,0,1,NA,37.321233,-120.65635400000001,0,20.45,0,0,Offer E,27808,0,0,0,0,1,1,0.0,43.82,0.0,20.45,0,0,95301
2829,1,1,0,0,8,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.7,560.85,1,80,22,14.89,3068,1,Ballico,0,1,Cable,37.4695,-120.672724,0,72.488,0,0,None,809,0,3,0,0,8,3,123.0,119.12,0.0,560.85,0,0,95303
2830,1,0,0,0,60,1,0,DSL,1,1,0,0,Two year,0,Electronic check,61.4,3638.25,0,24,26,30.92,6209,0,Big Oak Flat,1,1,Cable,37.818589,-120.25699499999999,0,61.4,0,0,Offer B,167,0,1,0,0,60,1,946.0,1855.2,0.0,3638.25,1,0,95305
2831,0,1,1,0,12,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,98.1,1060.2,1,67,30,30.63,2709,1,Catheys Valley,1,0,DSL,37.394411,-120.12726200000002,1,102.024,0,1,Offer D,986,0,2,1,0,12,5,318.0,367.56,49.06,1060.2,0,0,95306
2832,1,0,1,0,40,1,1,DSL,0,1,1,0,One year,0,Credit card (automatic),70.75,2921.75,0,33,22,23.74,5507,0,Ceres,0,1,Cable,37.553469,-120.952825,1,70.75,0,0,Offer B,32881,1,1,0,0,40,1,0.0,949.6,0.0,2921.75,0,1,95307
2833,0,0,0,0,66,1,0,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),61.15,4017.45,0,25,30,21.37,5133,0,Columbia,1,0,DSL,38.085839,-120.37855,0,61.15,0,0,None,2144,0,0,0,0,66,2,1205.0,1410.42,0.0,4017.45,1,0,95310
2834,1,0,1,1,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.25,854.9,0,57,0,9.33,4439,0,Coulterville,0,1,NA,37.722127,-120.110174,1,20.25,2,4,Offer B,2271,0,0,1,0,42,0,0.0,391.86,0.0,854.9,0,0,95311
2835,0,1,0,0,66,1,1,DSL,1,1,0,0,One year,1,Credit card (automatic),63.85,4174.35,0,72,5,36.48,4657,0,Cressey,0,0,Cable,37.420273,-120.66526999999999,0,63.85,0,0,Offer A,55,1,0,0,0,66,0,20.87,2407.68,0.0,4174.35,0,1,95312
2836,1,0,0,0,49,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,98.7,4920.55,0,56,27,45.46,6148,0,Crows Landing,0,1,Fiber Optic,37.435664,-121.04905600000001,0,98.7,0,0,Offer B,1508,0,0,0,1,49,1,0.0,2227.54,0.0,4920.55,0,1,95313
2837,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.5,20.5,1,24,0,26.12,3820,1,Delhi,0,0,NA,37.422961,-120.76549299999999,0,20.5,0,0,Offer E,10159,0,0,0,0,1,2,0.0,26.12,0.0,20.5,1,0,95315
2838,0,0,0,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.0,810.3,0,23,0,10.09,5913,0,Denair,0,0,NA,37.524721,-120.757977,0,20.0,0,0,Offer B,5513,0,1,0,0,41,2,0.0,413.69,0.0,810.3,1,0,95316
2839,0,0,1,1,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.3,772.4,0,34,0,21.28,4180,0,El Nido,0,0,NA,37.127386,-120.506422,1,19.3,1,1,Offer B,808,0,1,1,0,41,2,0.0,872.48,0.0,772.4,0,0,95317
2840,0,0,1,1,23,1,0,Fiber optic,1,1,0,0,Month-to-month,0,Mailed check,84.4,1936.85,0,19,82,27.24,2177,0,El Portal,0,0,Fiber Optic,37.654551,-119.822984,1,84.4,2,5,None,579,1,0,1,0,23,1,0.0,626.52,0.0,1936.85,1,1,95318
2841,1,0,0,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,25.1,79.8,0,28,69,0.0,2013,0,Escalon,0,1,Fiber Optic,37.818543,-121.00690700000001,0,25.1,0,0,Offer E,11474,0,0,0,0,3,0,0.0,0.0,0.0,79.8,1,1,95320
2842,0,0,0,0,4,0,No phone service,DSL,1,0,0,1,Month-to-month,0,Mailed check,48.25,202.25,0,19,30,0.0,2682,0,Groveland,1,0,Fiber Optic,37.902968,-119.66754399999999,0,48.25,0,0,Offer E,3680,1,0,0,1,4,0,61.0,0.0,0.0,202.25,1,0,95321
2843,0,0,1,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.85,1070.5,0,27,0,3.41,5432,0,Gustine,0,0,NA,37.147197999999996,-121.12016100000001,1,19.85,1,1,Offer B,7872,0,0,1,0,52,0,0.0,177.32,0.0,1070.5,1,0,95322
2844,0,1,1,0,4,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,99.6,347.65,1,68,22,18.91,4708,1,Hickman,0,0,Cable,37.605926000000004,-120.69955,1,103.584,0,1,None,1055,0,1,1,0,4,2,76.0,75.64,25.79,347.65,0,0,95323
2845,0,0,0,0,11,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,94.2,999.9,0,54,4,9.52,2405,0,Hilmar,1,0,Cable,37.394535999999995,-120.89074699999999,0,94.2,0,0,None,7177,1,0,0,1,11,0,40.0,104.72,0.0,999.9,0,0,95324
2846,0,0,1,0,2,1,0,DSL,1,0,0,1,Month-to-month,1,Mailed check,62.15,113.1,0,59,24,48.39,5766,0,Hornitos,0,0,Fiber Optic,37.479926,-120.230424,1,62.15,0,6,Offer E,128,0,0,1,1,2,2,27.0,96.78,0.0,113.1,0,0,95325
2847,0,0,1,0,26,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),79.3,2015.8,0,50,10,37.6,5168,0,Hughson,0,0,Fiber Optic,37.5923,-120.85328799999999,1,79.3,0,5,None,6822,0,0,1,0,26,0,20.16,977.6,0.0,2015.8,0,1,95326
2848,1,0,1,1,24,1,0,DSL,1,0,0,0,One year,1,Credit card (automatic),56.25,1454.25,0,33,53,2.31,3607,0,Jamestown,1,1,Cable,37.84771,-120.486589,1,56.25,3,7,None,9559,0,1,1,0,24,1,771.0,55.44,0.0,1454.25,0,0,95327
2849,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.3,246.7,0,26,0,32.32,4177,0,Keyes,0,0,NA,37.555631,-120.911653,0,20.3,0,0,None,2130,0,0,0,0,12,2,0.0,387.84,0.0,246.7,1,0,95328
2850,1,1,1,0,60,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.0,6017.9,0,69,5,10.4,4763,0,La Grange,0,1,DSL,37.666587,-120.41151699999999,1,99.0,0,5,Offer B,1749,1,0,1,0,60,2,0.0,624.0,0.0,6017.9,0,1,95329
2851,0,0,1,1,64,1,1,DSL,1,1,1,1,Two year,1,Mailed check,90.6,5817.45,0,44,19,37.0,5240,0,Lathrop,1,0,Fiber Optic,37.808209999999995,-121.308401,1,90.6,1,3,None,10834,1,0,1,1,64,0,0.0,2368.0,0.0,5817.45,0,1,95330
2852,1,0,1,0,66,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),85.9,5595.3,0,42,10,7.61,5137,0,Le Grand,1,1,DSL,37.249377,-120.249581,1,85.9,0,2,None,3256,1,0,1,1,66,0,560.0,502.2600000000001,0.0,5595.3,0,0,95333
2853,0,0,0,0,60,1,1,Fiber optic,0,0,0,0,One year,1,Bank transfer (automatic),79.2,4765,0,24,48,15.29,5687,0,Livingston,1,0,Fiber Optic,37.361987,-120.74839399999999,0,79.2,0,0,None,12672,0,0,0,0,60,1,0.0,917.4,0.0,4765.0,1,1,95334
2854,1,0,1,1,17,1,1,DSL,1,0,1,0,One year,1,Bank transfer (automatic),70.35,1201.65,0,36,76,33.24,2704,0,Long Barn,1,1,DSL,38.109125,-120.078597,1,70.35,3,5,None,683,0,0,1,0,17,3,0.0,565.08,0.0,1201.65,0,1,95335
2855,1,0,1,1,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.35,867.3,0,63,0,34.33,3433,0,Manteca,0,1,NA,37.830267,-121.20101799999999,1,19.35,2,10,None,36738,0,0,1,0,42,0,0.0,1441.86,0.0,867.3,0,0,95336
2856,1,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.15,50.15,0,42,2,39.87,3043,0,Manteca,0,1,DSL,37.750822,-121.238423,0,50.15,0,0,Offer E,19867,0,1,0,0,1,2,0.0,39.87,0.0,50.15,0,1,95337
2857,0,0,1,1,47,1,0,DSL,0,1,0,1,Two year,0,Bank transfer (automatic),63.8,3007.25,0,32,57,30.06,5144,0,Mariposa,0,0,DSL,37.526790999999996,-119.99436999999999,1,63.8,3,0,None,10226,1,0,0,1,47,1,171.41,1412.82,0.0,3007.25,0,1,95338
2858,0,0,1,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.55,252.75,0,27,0,10.42,4907,0,Merced,0,0,NA,37.255637,-120.49353700000002,1,20.55,0,2,None,59289,0,1,1,0,10,4,0.0,104.2,0.0,252.75,1,0,95340
2859,1,1,1,0,70,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),88.55,6306.5,0,69,8,40.94,4097,0,Midpines,1,1,Fiber Optic,37.581496,-119.97276200000002,1,88.55,0,4,None,433,1,0,1,0,70,0,505.0,2865.8,0.0,6306.5,0,0,95345
2860,1,1,0,0,67,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),101.4,6841.05,0,76,19,38.85,5269,0,Mi Wuk Village,1,1,Fiber Optic,38.121601,-120.13391499999999,0,101.4,0,0,None,1278,0,0,0,0,67,2,1300.0,2602.9500000000007,0.0,6841.05,0,0,95346
2861,0,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,81.95,81.95,1,44,18,44.94,5622,1,Merced,0,0,DSL,37.40122,-120.514191,0,85.22800000000002,0,0,Offer E,23100,0,4,0,1,1,4,0.0,44.94,0.0,81.95,0,0,95348
2862,1,0,1,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.35,451.1,1,39,31,14.75,4292,1,Modesto,0,1,Cable,37.671806,-121.007575,1,72.124,0,1,Offer E,52872,0,0,1,0,7,0,140.0,103.25,0.0,451.1,0,0,95350
2863,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.6,44.6,0,45,2,45.28,4864,0,Modesto,0,1,DSL,37.621458000000004,-121.012295,0,44.6,0,0,None,47536,0,0,0,0,1,1,0.0,45.28,0.0,44.6,0,1,95351
2864,1,0,0,0,4,1,0,DSL,0,1,1,0,Month-to-month,1,Bank transfer (automatic),63.75,226.2,0,53,11,3.03,2624,0,Modesto,0,1,Fiber Optic,37.639029,-120.964772,0,63.75,0,0,None,27135,1,0,0,0,4,0,25.0,12.12,0.0,226.2,0,0,95354
2865,0,0,1,1,66,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),109.25,7082.5,0,61,25,20.11,5865,0,Modesto,1,0,Cable,37.672906,-120.94659399999999,1,109.25,2,2,None,47613,0,0,1,1,66,1,0.0,1327.26,0.0,7082.5,0,1,95355
2866,0,0,0,0,12,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,84.6,1017.35,0,31,25,2.57,4807,0,Modesto,0,0,Fiber Optic,37.716186,-121.02583600000001,0,84.6,0,0,None,26055,0,1,0,1,12,1,254.0,30.84,0.0,1017.35,0,0,95356
2867,0,0,0,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.45,527.35,0,25,0,5.98,4690,0,Modesto,0,0,NA,37.670526,-120.877572,0,20.45,0,0,None,13343,0,0,0,0,24,0,0.0,143.52,0.0,527.35,1,0,95357
2868,1,0,0,0,26,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,85.75,2146.5,0,48,13,40.35,3178,0,Modesto,0,1,DSL,37.612612,-121.10856799999999,0,85.75,0,0,None,30668,0,0,0,0,26,0,27.9,1049.1,0.0,2146.5,0,1,95358
2869,0,0,0,0,6,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,91.1,455.3,1,53,26,11.81,2266,1,Newman,0,0,Cable,37.343846,-121.039391,0,94.744,0,0,None,8504,0,2,0,1,6,1,118.0,70.86,0.0,455.3,0,0,95360
2870,1,0,1,0,57,1,1,Fiber optic,0,0,1,1,Two year,0,Electronic check,107.95,5969.85,0,31,29,16.78,4687,0,Oakdale,1,1,Fiber Optic,37.785033,-120.776141,1,107.95,0,2,None,25384,1,0,1,1,57,1,0.0,956.46,0.0,5969.85,0,1,95361
2871,1,0,1,0,14,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.1,1235.55,1,20,46,7.26,2177,1,Patterson,0,1,Fiber Optic,37.410236,-121.32033700000001,1,89.544,0,1,Offer D,15536,0,2,1,0,14,2,568.0,101.64,0.0,1235.55,1,0,95363
2872,0,0,1,1,42,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,22.95,1014.25,0,47,0,13.95,4650,0,Pinecrest,0,0,NA,38.224869,-119.755729,1,22.95,3,1,None,235,0,1,1,0,42,2,0.0,585.9,0.0,1014.25,0,0,95364
2873,1,0,0,0,25,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),94.7,2362.1,1,41,9,34.88,5641,1,Planada,0,1,Cable,37.329725,-120.306399,0,98.488,0,0,None,4150,0,3,0,1,25,2,213.0,872.0000000000001,0.0,2362.1,0,0,95365
2874,0,0,1,0,64,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.45,1225.65,0,25,0,14.78,5113,0,Ripon,0,0,NA,37.750778000000004,-121.13238,1,19.45,0,4,None,12646,0,0,1,0,64,0,0.0,945.92,0.0,1225.65,1,0,95366
2875,1,0,1,0,22,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.1,1873.7,1,40,19,16.2,5248,1,Riverbank,0,1,Cable,37.734971,-120.95427099999999,1,88.50399999999998,0,1,Offer D,16525,0,3,1,1,22,3,0.0,356.4,0.0,1873.7,0,1,95367
2876,1,0,0,0,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),19.7,386.5,0,62,0,26.54,4431,0,Salida,0,1,NA,37.713152,-121.08738999999998,0,19.7,0,0,None,12466,0,0,0,0,19,0,0.0,504.26,0.0,386.5,0,0,95368
2877,0,0,1,1,61,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.15,6010.05,1,63,8,49.33,5612,1,Snelling,0,0,Cable,37.521708000000004,-120.42684299999999,1,103.116,0,1,None,1158,0,0,1,1,61,0,48.08,3009.13,0.0,6010.05,0,1,95369
2878,1,0,1,0,22,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),87.0,1850.65,0,56,18,48.68,5233,0,Sonora,1,1,Fiber Optic,37.982715999999996,-120.343732,1,87.0,0,9,None,25340,0,0,1,0,22,2,0.0,1070.96,0.0,1850.65,0,1,95370
2879,1,1,1,0,70,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,102.95,7101.5,1,69,22,17.45,5005,1,Soulsbyville,1,1,DSL,37.990574,-120.261821,1,107.068,0,1,None,1519,0,4,1,0,70,3,1562.0,1221.5,15.24,7101.5,0,0,95372
2880,1,0,0,0,12,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),79.95,1043.4,0,23,41,40.06,2968,0,Stevinson,0,1,DSL,37.316807,-120.855753,0,79.95,0,0,None,1960,0,0,0,1,12,0,428.0,480.72,0.0,1043.4,1,0,95374
2881,0,0,1,0,31,1,0,DSL,1,0,0,1,One year,1,Electronic check,64.0,1910.75,0,55,15,28.8,5191,0,Tracy,0,0,Fiber Optic,37.680968,-121.446049,1,64.0,0,9,None,69801,1,0,1,1,31,0,0.0,892.8000000000002,0.0,1910.75,0,1,95376
2882,0,0,0,0,11,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,64.9,716.1,0,42,17,13.56,2775,0,Tuolumne,0,0,DSL,37.939768,-120.188002,0,64.9,0,0,Offer D,3979,0,0,0,1,11,0,122.0,149.16,0.0,716.1,0,0,95379
2883,1,0,1,1,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.75,1686.15,0,36,0,26.83,5434,0,Turlock,0,1,NA,37.474396,-120.87591699999999,1,25.75,1,10,None,40545,0,0,1,0,68,0,0.0,1824.44,0.0,1686.15,0,0,95380
2884,0,1,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),90.15,6716.45,0,78,16,9.88,4606,0,Turlock,1,0,DSL,37.529656,-120.85435700000001,1,90.15,1,2,None,24708,1,0,1,0,72,0,1075.0,711.36,0.0,6716.45,0,0,95382
2885,1,1,0,0,67,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),116.1,7839.85,0,68,29,44.56,5896,0,Twain Harte,1,1,Cable,38.107440999999994,-120.230625,0,116.1,0,0,None,4848,1,0,0,0,67,0,0.0,2985.52,0.0,7839.85,0,1,95383
2886,0,0,0,0,60,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),104.95,6236.75,0,30,48,22.88,5926,0,Vernalis,1,0,Fiber Optic,37.609095,-121.26338100000001,0,104.95,0,0,None,274,1,0,0,1,60,1,0.0,1372.8,0.0,6236.75,0,1,95385
2887,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.05,45.05,1,31,29,13.84,2644,1,Waterford,0,1,Cable,37.669515999999994,-120.62696399999999,0,46.852,0,0,None,8308,0,1,0,0,1,2,0.0,13.84,0.0,45.05,0,0,95386
2888,0,1,0,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.0,71,1,80,6,28.64,5345,1,Escondido,0,0,DSL,33.141265000000004,-116.967221,0,73.84,0,0,None,48690,0,0,0,0,1,3,0.0,28.64,0.0,71.0,0,1,92027
2889,1,0,1,1,58,0,No phone service,DSL,1,1,1,0,One year,0,Mailed check,50.0,2919.85,0,21,52,0.0,4704,0,Winton,1,1,Cable,37.421299,-120.59958700000001,1,50.0,3,9,None,11463,0,0,1,0,58,0,0.0,0.0,0.0,2919.85,1,1,95388
2890,0,1,1,1,47,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),70.55,3309.25,1,73,29,26.95,4457,1,Escondido,0,0,Fiber Optic,33.141265000000004,-116.967221,1,73.372,0,1,None,48690,0,0,1,0,47,0,960.0,1266.65,26.99,3309.25,0,0,92027
2891,0,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.7,79.7,1,39,29,33.88,2066,1,Santa Rosa,0,0,Cable,38.460516999999996,-122.79033500000001,0,82.88799999999999,0,0,None,36125,0,1,0,1,1,2,0.0,33.88,0.0,79.7,0,0,95401
2892,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.45,20.45,0,32,0,39.61,2664,0,Santa Rosa,0,1,NA,38.488431,-122.752839,0,20.45,0,0,None,40270,0,0,0,0,1,1,0.0,39.61,0.0,20.45,0,0,95403
2893,1,0,0,0,22,1,1,DSL,1,1,0,0,Month-to-month,0,Electronic check,59.0,1254.7,1,46,19,49.43,2195,1,Santa Rosa,0,1,Cable,38.526941,-122.709096,0,61.36,0,0,Offer D,35057,0,1,0,0,22,5,238.0,1087.46,0.0,1254.7,0,0,95404
2894,0,0,0,0,48,1,0,DSL,1,0,0,0,One year,1,Credit card (automatic),60.35,2896.4,1,51,14,33.91,2681,1,Santa Rosa,1,0,Fiber Optic,38.439696000000005,-122.66881699999999,0,62.763999999999996,0,0,None,22250,1,0,0,0,48,4,0.0,1627.6799999999996,0.0,2896.4,0,1,95405
2895,0,0,1,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.85,717.5,0,54,0,15.51,5707,0,Santa Rosa,0,0,NA,38.394090999999996,-122.739814,1,19.85,0,8,None,30876,0,0,1,0,37,3,0.0,573.87,0.0,717.5,0,0,95407
2896,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,19.95,253.8,0,34,0,7.33,2252,0,Santa Rosa,0,1,NA,38.468893,-122.58053899999999,0,19.95,0,0,Offer D,25718,0,0,0,0,13,0,0.0,95.29,0.0,253.8,0,0,95409
2897,1,0,0,0,43,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),26.45,1110.05,0,39,0,28.9,3881,0,Albion,0,1,NA,39.225694,-123.717354,0,26.45,0,0,None,1054,0,1,0,0,43,2,0.0,1242.7,0.0,1110.05,0,0,95410
2898,0,0,0,0,6,0,No phone service,DSL,1,1,1,1,Two year,1,Mailed check,63.4,348.8,0,21,52,0.0,3909,0,Annapolis,1,0,Fiber Optic,38.731055,-123.316553,0,63.4,0,0,None,747,1,0,0,1,6,0,18.14,0.0,0.0,348.8,1,1,95412
2899,1,0,0,0,71,0,No phone service,DSL,1,1,1,0,Two year,0,Bank transfer (automatic),53.95,3888.65,0,46,20,0.0,4094,0,Boonville,1,1,Cable,39.025867,-123.38154399999999,0,53.95,0,0,None,1374,1,0,0,0,71,0,0.0,0.0,0.0,3888.65,0,1,95415
2900,0,1,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.25,69.25,1,73,9,37.3,4568,1,Branscomb,0,0,Fiber Optic,39.710591,-123.682799,1,72.02,0,1,None,176,0,3,1,0,1,1,0.0,37.3,0.0,69.25,0,0,95417
2901,0,0,1,1,72,1,1,Fiber optic,1,1,1,0,Two year,1,Electronic check,95.1,6843.15,0,39,19,18.74,5584,0,Caspar,0,0,Fiber Optic,39.361283,-123.784599,1,95.1,2,8,None,333,0,0,1,0,72,1,0.0,1349.28,0.0,6843.15,0,1,95420
2902,0,1,0,0,6,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,74.1,450.9,0,65,20,12.67,4716,0,Cazadero,0,0,DSL,38.578807,-123.19338,0,74.1,0,0,None,1575,0,0,0,0,6,0,9.02,76.02,0.0,450.9,0,1,95421
2903,1,0,1,1,12,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Mailed check,35.5,432.25,0,19,73,0.0,2562,0,Clearlake,0,1,DSL,38.965804,-122.63177900000001,1,35.5,3,7,Offer D,13485,1,0,1,0,12,2,0.0,0.0,0.0,432.25,1,1,95422
2904,1,0,0,0,25,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.95,1767.35,1,52,20,24.91,4881,1,Clearlake Oaks,0,1,Cable,39.07116,-122.598542,0,73.78800000000003,0,0,None,3684,0,1,0,0,25,2,353.0,622.75,0.0,1767.35,0,0,95423
2905,0,0,1,0,21,1,0,Fiber optic,0,0,0,0,One year,0,Electronic check,79.2,1742.45,0,49,20,14.51,4900,0,Cloverdale,1,0,Fiber Optic,38.801936,-122.93893500000001,1,79.2,0,7,Offer D,9210,1,0,1,0,21,0,0.0,304.71,0.0,1742.45,0,1,95425
2906,0,0,1,1,6,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,48.8,297.35,0,39,10,49.45,4538,0,Cobb,0,0,Fiber Optic,38.838088,-122.73203000000001,1,48.8,2,3,None,1591,1,0,1,0,6,1,2.97,296.7000000000001,0.0,297.35,0,1,95426
2907,1,0,1,0,20,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,89.0,1820.45,1,35,6,18.05,4594,1,Comptche,0,1,DSL,39.239818,-123.565432,1,92.56,0,1,Offer D,371,0,2,1,1,20,2,0.0,361.0,0.0,1820.45,0,1,95427
2908,1,0,1,0,18,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,99.4,1742.95,1,51,18,11.3,2421,1,Covelo,0,1,Cable,39.83307,-123.17876499999998,1,103.376,0,1,None,2296,0,0,1,1,18,2,314.0,203.4,0.0,1742.95,0,0,95428
2909,0,0,0,0,43,1,0,DSL,0,1,0,0,One year,0,Electronic check,55.45,2444.25,0,38,19,1.6,3350,0,Dos Rios,0,0,Cable,39.756049,-123.358701,0,55.45,0,0,None,91,1,0,0,0,43,1,464.0,68.8,0.0,2444.25,0,0,95429
2910,0,0,1,1,35,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.4,949.8,0,53,0,32.75,5070,0,Duncans Mills,0,0,NA,38.445603000000006,-123.06375600000001,1,25.4,1,9,None,187,0,0,1,0,35,0,0.0,1146.25,0.0,949.8,0,0,95430
2911,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),73.5,73.5,1,50,2,3.84,4378,1,Eldridge,1,0,DSL,38.348884000000005,-122.51698999999999,0,76.44,0,0,None,363,0,2,0,0,1,1,0.0,3.84,0.0,73.5,0,1,95431
2912,1,1,1,0,32,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,93.5,2970.8,0,78,3,43.54,5804,0,Elk,1,1,Cable,39.108252,-123.645121,1,93.5,0,9,Offer C,383,0,0,1,0,32,0,89.0,1393.28,0.0,2970.8,0,0,95432
2913,1,0,0,0,52,0,No phone service,DSL,1,1,1,1,Two year,0,Credit card (automatic),63.9,3334.95,0,57,18,0.0,5380,0,Forestville,1,1,Cable,38.499302,-122.92443999999999,0,63.9,0,0,None,6216,1,0,0,1,52,0,0.0,0.0,0.0,3334.95,0,1,95436
2914,1,0,0,0,32,1,0,DSL,0,0,1,1,One year,1,Bank transfer (automatic),64.85,2010.95,0,43,12,15.52,4895,0,Fort Bragg,0,1,Fiber Optic,39.455555,-123.68397900000001,0,64.85,0,0,None,14417,0,0,0,1,32,1,0.0,496.64,0.0,2010.95,0,1,95437
2915,0,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),63.8,4684.3,0,61,22,0.0,6107,0,Fulton,1,0,Fiber Optic,38.493888,-122.77714099999999,1,63.8,3,8,None,476,1,0,1,1,72,2,1031.0,0.0,0.0,4684.3,0,0,95439
2916,1,0,0,0,51,0,No phone service,DSL,1,0,0,1,Month-to-month,1,Credit card (automatic),44.45,2181.55,0,31,2,0.0,6087,0,Geyserville,0,1,Fiber Optic,38.731771,-123.064272,0,44.45,0,0,None,2349,1,0,0,1,51,0,0.0,0.0,0.0,2181.55,0,1,95441
2917,1,0,1,1,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.95,1303.25,0,47,0,19.75,6492,0,Glen Ellen,0,1,NA,38.368744,-122.52264199999999,1,19.95,3,4,Offer A,4101,0,0,1,0,68,1,0.0,1343.0,0.0,1303.25,0,0,95442
2918,1,1,1,0,8,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Mailed check,43.35,371.4,0,67,27,0.0,2560,0,Glenhaven,1,1,Cable,39.045246,-122.743181,1,43.35,0,1,None,175,0,0,1,0,8,0,10.03,0.0,0.0,371.4,0,1,95443
2919,1,0,1,0,49,0,No phone service,DSL,0,1,1,1,Two year,0,Credit card (automatic),49.65,2409.9,0,22,27,0.0,4283,0,Graton,0,1,DSL,38.434362,-122.86891000000001,1,49.65,0,8,None,390,0,0,1,1,49,1,0.0,0.0,0.0,2409.9,1,1,95444
2920,0,0,1,0,72,1,0,DSL,1,1,1,1,Two year,0,Mailed check,85.1,6155.4,0,24,41,20.54,4147,0,Gualala,1,0,Cable,38.848082,-123.50608000000001,1,85.1,0,7,Offer A,1916,1,0,1,1,72,0,2524.0,1478.88,0.0,6155.4,1,0,95445
2921,1,0,0,0,9,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.5,829.1,1,45,11,19.22,5007,1,Guerneville,0,1,Cable,38.52576,-123.013347,0,99.32,0,0,None,4913,0,3,0,1,9,2,9.12,172.98,0.0,829.1,0,1,95446
2922,0,0,1,0,28,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Mailed check,92.35,2602.9,1,47,22,37.66,2990,1,Healdsburg,0,0,Cable,38.618347,-122.908422,1,96.044,0,1,None,17979,0,2,1,1,28,2,573.0,1054.48,0.0,2602.9,0,0,95448
2923,1,0,0,0,54,1,0,Fiber optic,1,0,1,0,Month-to-month,0,Mailed check,89.8,4667,0,55,24,27.17,4980,0,Hopland,1,1,Fiber Optic,38.937059999999995,-123.11811100000001,0,89.8,0,0,None,1373,0,0,0,0,54,0,0.0,1467.18,0.0,4667.0,0,1,95449
2924,1,0,0,0,11,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.55,824.75,1,20,45,5.4,4601,1,Jenner,0,1,DSL,38.505995,-123.18701899999999,0,77.532,0,0,None,438,0,2,0,0,11,2,0.0,59.40000000000001,0.0,824.75,1,1,95450
2925,0,0,1,1,50,1,0,Fiber optic,0,0,1,1,One year,0,Mailed check,103.05,5153.5,0,41,27,47.48,5905,0,Kelseyville,1,0,Fiber Optic,38.93496,-122.792243,1,103.05,3,7,None,9902,1,0,1,1,50,0,1391.0,2374.0,0.0,5153.5,0,0,95451
2926,0,0,1,0,69,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,116.0,8182.85,0,55,27,38.52,4216,0,Kenwood,1,0,Fiber Optic,38.419525,-122.52158500000002,1,116.0,0,3,Offer A,1653,1,0,1,1,69,0,2209.0,2657.88,0.0,8182.85,0,0,95452
2927,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.9,69.9,0,46,14,9.36,3358,0,Lakeport,0,1,Cable,39.080469,-122.955176,0,69.9,0,0,None,11180,0,1,0,0,1,4,0.0,9.36,0.0,69.9,0,1,95453
2928,1,0,1,1,68,1,0,Fiber optic,1,1,0,1,Two year,0,Bank transfer (automatic),95.1,6683.4,0,31,18,9.29,5748,0,Laytonville,0,1,Fiber Optic,39.806141,-123.531098,1,95.1,2,3,Offer A,2706,1,0,1,1,68,1,120.3,631.7199999999998,0.0,6683.4,0,1,95454
2929,1,0,0,1,40,0,No phone service,DSL,1,1,0,0,One year,0,Mailed check,40.25,1564.05,0,62,57,0.0,4288,0,Little River,0,1,Fiber Optic,39.245911,-123.77214,0,40.25,3,0,None,882,1,0,0,0,40,0,89.15,0.0,0.0,1564.05,0,1,95456
2930,1,0,1,1,31,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.75,755.6,0,26,0,7.03,5472,0,Lower Lake,0,1,NA,38.925545,-122.54908300000001,1,25.75,3,7,None,2644,0,0,1,0,31,0,0.0,217.93,0.0,755.6,1,0,95457
2931,0,1,0,1,33,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),105.35,3465.05,0,73,19,12.75,4738,0,Lucerne,1,0,Fiber Optic,39.141934,-122.770679,0,105.35,2,0,Offer C,3002,0,0,0,0,33,0,658.0,420.75,0.0,3465.05,0,0,95458
2932,1,1,1,0,55,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,113.6,6292.7,0,72,21,12.91,5754,0,Manchester,1,1,DSL,38.966713,-123.58641200000001,1,113.6,0,7,Offer B,586,1,0,1,0,55,0,0.0,710.05,0.0,6292.7,0,1,95459
2933,1,0,1,1,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.0,1664.3,0,60,0,2.71,5440,0,Mendocino,0,1,NA,39.305545,-123.743697,1,24.0,1,8,Offer A,2229,0,0,1,0,68,2,0.0,184.28,0.0,1664.3,0,0,95460
2934,0,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.4,198.1,0,48,0,8.25,3713,0,Middletown,0,0,NA,38.787446,-122.58675,1,19.4,1,0,Offer D,7789,0,0,0,0,12,0,0.0,99.0,0.0,198.1,0,0,95461
2935,1,0,1,0,71,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),86.1,6045.9,0,39,6,5.51,6286,0,Monte Rio,1,1,DSL,38.471049,-123.015549,1,86.1,0,7,Offer A,1537,1,0,1,1,71,1,36.28,391.21,0.0,6045.9,0,1,95462
2936,1,0,0,0,40,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Mailed check,102.65,4108.15,0,42,29,32.78,3655,0,Navarro,1,1,Fiber Optic,39.182916,-123.552571,0,102.65,0,0,None,148,0,1,0,1,40,1,1191.0,1311.2,0.0,4108.15,0,0,95463
2937,0,0,1,1,64,1,1,Fiber optic,0,1,0,1,One year,1,Electronic check,92.85,5980.75,0,21,69,37.47,5206,0,Nice,1,0,Fiber Optic,39.12334,-122.83819799999999,1,92.85,3,8,None,2223,0,0,1,1,64,0,0.0,2398.08,0.0,5980.75,1,1,95464
2938,1,0,1,0,53,1,1,Fiber optic,0,1,0,1,One year,0,Bank transfer (automatic),97.75,5043.2,0,44,17,32.94,4488,0,Occidental,0,1,Fiber Optic,38.415003000000006,-122.998726,1,97.75,0,6,None,1880,1,0,1,1,53,0,0.0,1745.82,0.0,5043.2,0,1,95465
2939,1,1,0,0,12,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,83.8,1029.75,1,65,8,28.63,5565,1,Philo,1,1,Fiber Optic,39.094102,-123.500853,0,87.152,0,0,Offer D,1113,1,3,0,0,12,4,82.0,343.56,44.58,1029.75,0,0,95466
2940,1,1,0,0,53,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,54.45,2854.55,1,73,28,0.0,6280,1,Point Arena,1,1,DSL,38.911299,-123.60958799999999,0,56.62800000000001,0,0,None,1352,0,0,0,0,53,0,799.0,0.0,20.16,2854.55,0,0,95468
2941,1,0,1,0,72,1,1,Fiber optic,1,1,1,0,Two year,1,Credit card (automatic),97.95,7114.25,0,43,3,38.3,4256,0,Potter Valley,1,1,Fiber Optic,39.408634,-123.04551599999999,1,97.95,0,1,Offer A,1884,0,0,1,0,72,1,213.0,2757.6,0.0,7114.25,0,0,95469
2942,1,0,0,0,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,19.95,907.05,0,51,0,13.42,4006,0,Redwood Valley,0,1,NA,39.298065,-123.25211000000002,0,19.95,0,0,None,5995,0,0,0,0,46,0,0.0,617.32,0.0,907.05,0,0,95470
2943,1,0,0,0,40,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.6,973.95,0,27,0,27.47,2601,0,Rio Nido,0,1,NA,38.522328,-122.97932,0,24.6,0,0,None,298,0,0,0,0,40,0,0.0,1098.8,0.0,973.95,1,0,95471
2944,1,0,0,0,12,0,No phone service,DSL,1,1,1,0,Month-to-month,1,Bank transfer (automatic),50.95,605.75,0,45,9,0.0,2716,0,Sebastopol,0,1,Cable,38.398815,-122.861923,0,50.95,0,0,Offer D,31266,1,0,0,0,12,0,0.0,0.0,0.0,605.75,0,1,95472
2945,1,0,0,0,9,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,75.6,661.55,0,58,6,21.11,4990,0,Sonoma,0,1,Fiber Optic,38.25485,-122.461799,0,75.6,0,0,None,34314,0,0,0,0,9,3,0.0,189.99,0.0,661.55,0,1,95476
2946,0,0,1,1,51,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,80.75,4116.9,0,40,27,29.56,6032,0,Ukiah,0,0,Fiber Optic,39.134075,-123.23422,1,80.75,2,9,Offer B,30988,1,1,1,0,51,1,111.16,1507.56,0.0,4116.9,0,1,95482
2947,1,0,1,1,49,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),90.4,4494.65,0,62,20,11.74,5804,0,Upper Lake,1,1,Cable,39.220368,-122.907693,1,90.4,3,10,Offer B,2344,0,0,1,0,49,0,89.89,575.26,0.0,4494.65,0,1,95485
2948,1,1,1,0,41,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.8,4259.3,1,78,16,22.56,4726,1,Westport,1,1,DSL,39.724433000000005,-123.767578,1,103.792,0,0,None,309,0,4,0,0,41,4,681.0,924.96,8.88,4259.3,0,0,95488
2949,0,0,0,0,56,1,0,DSL,1,0,0,0,One year,1,Credit card (automatic),60.25,3282.75,0,32,22,30.86,4835,0,Willits,1,0,Fiber Optic,39.492046,-123.375818,0,60.25,0,0,Offer B,13472,1,0,0,0,56,1,722.0,1728.16,0.0,3282.75,0,0,95490
2950,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.2,55.7,0,29,0,46.53,4267,0,Windsor,0,1,NA,38.527297,-122.81004399999999,0,20.2,0,0,None,23701,0,2,0,0,4,2,0.0,186.12,0.0,55.7,1,0,95492
2951,1,0,1,0,20,1,0,DSL,1,0,0,1,One year,1,Mailed check,64.15,1274.45,0,45,18,33.78,5969,0,Witter Springs,0,1,Cable,39.222322999999996,-122.98548799999999,1,64.15,0,3,Offer D,240,1,0,1,1,20,1,22.94,675.6,0.0,1274.45,0,1,95493
2952,0,0,1,1,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.25,493.95,0,41,0,24.44,5158,0,Yorkville,0,0,NA,38.888351,-123.23964699999999,1,20.25,1,4,None,335,0,0,1,0,26,1,0.0,635.44,0.0,493.95,0,0,95494
2953,0,0,1,1,20,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),105.85,2239.65,1,57,18,28.79,4223,1,The Sea Ranch,1,0,Cable,38.696659000000004,-123.43686100000001,1,110.084,0,3,None,752,0,4,1,1,20,4,403.0,575.8,0.0,2239.65,0,0,95497
2954,0,0,0,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,75.45,480.75,1,35,16,18.1,2872,1,Eureka,0,0,Fiber Optic,40.796621,-124.15428,0,78.468,0,0,None,23224,0,0,0,0,7,0,77.0,126.70000000000002,0.0,480.75,0,0,95501
2955,1,0,0,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.85,635.6,1,60,25,15.51,3506,1,Eureka,0,1,DSL,40.737431,-124.108897,0,97.604,0,0,None,23570,0,2,0,1,7,3,159.0,108.57,0.0,635.6,0,0,95503
2956,1,0,0,0,51,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.0,5038.15,0,34,2,42.33,5787,0,Alderpoint,1,1,Cable,40.166028000000004,-123.584144,0,99.0,0,0,Offer B,261,0,2,0,1,51,2,0.0,2158.83,0.0,5038.15,0,1,95511
2957,0,0,0,0,4,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,80.3,324.2,0,26,51,38.74,3132,0,Blocksburg,0,0,Fiber Optic,40.309088,-123.668201,0,80.3,0,0,None,199,0,2,0,0,4,1,165.0,154.96,0.0,324.2,1,0,95514
2958,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.55,19.55,0,30,0,8.23,5537,0,Mckinleyville,0,0,NA,40.965011,-124.01525500000001,0,19.55,0,0,None,15921,0,0,0,0,1,2,0.0,8.23,0.0,19.55,0,0,95519
2959,1,0,1,1,27,1,1,Fiber optic,1,1,1,0,Month-to-month,0,Electronic check,100.75,2793.55,0,39,15,14.07,3160,0,Arcata,0,1,Fiber Optic,40.839958,-124.00375700000001,1,100.75,1,0,None,19596,1,0,0,0,27,2,0.0,379.89,0.0,2793.55,0,1,95521
2960,1,0,0,0,22,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,100.75,2095,1,51,19,35.93,4152,1,Bayside,0,1,Cable,40.825486,-124.049485,0,104.78,0,0,None,1689,0,1,0,1,22,3,398.0,790.46,0.0,2095.0,0,0,95524
2961,1,0,0,0,12,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,53.75,648.65,0,53,3,1.8,5385,0,Blue Lake,0,1,Fiber Optic,40.94338,-123.831799,0,53.75,0,0,Offer D,1584,1,0,0,0,12,1,19.0,21.6,0.0,648.65,0,0,95525
2962,0,0,1,1,3,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,31.0,95.05,1,43,21,0.0,5122,1,Bridgeville,0,0,Fiber Optic,40.372532,-123.525626,1,32.24,1,1,None,695,1,0,1,0,3,1,0.0,0.0,0.0,95.05,0,1,95526
2963,0,0,1,1,34,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),25.6,917.15,0,57,0,25.69,5854,0,Burnt Ranch,0,0,NA,40.854512,-123.450097,1,25.6,1,6,None,485,0,0,1,0,34,2,0.0,873.46,0.0,917.15,0,0,95527
2964,1,0,1,0,24,1,1,DSL,1,0,0,0,One year,1,Electronic check,58.35,1346.9,0,50,4,34.01,5428,0,Carlotta,0,1,Fiber Optic,40.497283,-123.93037,1,58.35,0,5,None,1072,1,0,1,0,24,0,0.0,816.24,0.0,1346.9,0,1,95528
2965,1,0,0,0,51,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),80.0,4242.35,1,38,18,5.62,4769,1,Fallbrook,1,1,Fiber Optic,33.362575,-117.299644,0,83.2,0,0,None,42239,0,0,0,0,51,1,764.0,286.62,0.0,4242.35,0,0,92028
2966,0,1,0,0,14,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,46.35,672.7,0,71,5,0.0,2056,0,Ferndale,0,0,Fiber Optic,40.4785,-124.301372,0,46.35,0,0,None,2965,0,0,0,1,14,2,34.0,0.0,0.0,672.7,0,0,95536
2967,1,0,1,0,59,1,1,Fiber optic,1,1,1,1,Two year,0,Electronic check,113.75,6561.25,0,34,19,14.98,6251,0,Fields Landing,1,1,DSL,40.726949,-124.217378,1,113.75,0,9,Offer B,228,1,0,1,1,59,1,0.0,883.82,0.0,6561.25,0,1,95537
2968,1,0,0,0,3,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,90.4,268.45,0,22,73,31.48,5625,0,Fortuna,1,1,DSL,40.584990999999995,-124.121504,0,90.4,0,0,None,12241,0,0,0,1,3,1,196.0,94.44,0.0,268.45,1,0,95540
2969,0,0,1,1,65,1,1,Fiber optic,1,0,1,1,Two year,0,Electronic check,109.3,7337.55,0,22,47,13.25,6087,0,Garberville,1,0,Cable,40.057784000000005,-123.679461,1,109.3,2,4,Offer B,2423,1,0,1,1,65,0,3449.0,861.25,0.0,7337.55,1,0,95542
2970,1,1,0,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.25,331.9,1,68,19,2.27,3684,1,Gasquet,0,1,Cable,41.867908,-123.79414399999999,0,73.06,0,0,None,532,0,0,0,0,5,0,0.0,11.35,12.48,331.9,0,1,95543
2971,0,0,1,1,59,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),90.3,5194.05,0,50,24,47.05,4617,0,Honeydew,1,0,DSL,40.342928,-124.06332900000001,1,90.3,2,5,Offer B,82,1,0,1,1,59,0,124.66,2775.95,0.0,5194.05,0,1,95545
2972,1,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,1,Credit card (automatic),65.25,4478.85,0,24,51,0.0,6412,0,Hoopa,1,1,DSL,41.163637,-123.70484099999999,1,65.25,3,9,Offer A,3041,1,0,1,1,72,0,0.0,0.0,0.0,4478.85,1,1,95546
2973,0,0,1,1,62,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.15,6283.3,1,32,14,48.58,4120,1,Hydesville,1,0,Cable,40.557314,-124.08166200000001,1,104.156,0,1,None,1201,0,2,1,1,62,3,880.0,3011.96,0.0,6283.3,0,0,95547
2974,1,0,0,0,28,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Credit card (automatic),94.5,2659.4,1,52,29,35.52,5433,1,Klamath,0,1,Fiber Optic,41.572813000000004,-124.03501100000001,0,98.28,0,0,None,1215,0,2,0,1,28,3,771.0,994.56,0.0,2659.4,0,0,95548
2975,1,0,0,0,3,1,0,DSL,0,0,0,1,Month-to-month,0,Mailed check,60.65,196.9,0,43,11,22.49,2111,0,Kneeland,0,1,Fiber Optic,40.664483000000004,-123.865325,0,60.65,0,0,None,264,1,0,0,1,3,1,2.17,67.47,0.0,196.9,0,1,95549
2976,1,0,0,1,19,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),24.1,439.2,0,62,0,14.48,2378,0,Korbel,0,1,NA,40.7666,-123.80458,0,24.1,2,0,Offer D,155,0,0,0,0,19,2,0.0,275.12,0.0,439.2,0,0,95550
2977,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.5,19.5,0,54,0,8.02,3753,0,Loleta,0,1,NA,40.665952000000004,-124.240051,0,19.5,0,0,None,1447,0,0,0,0,1,0,0.0,8.02,0.0,19.5,0,0,95551
2978,1,0,0,0,24,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,85.95,2107.15,0,60,24,9.53,5421,0,Mad River,1,1,DSL,40.390301,-123.412327,0,85.95,0,0,None,265,1,0,0,0,24,2,0.0,228.72,0.0,2107.15,0,1,95552
2979,1,1,0,0,57,1,0,DSL,0,0,0,0,One year,1,Electronic check,53.5,3035.8,0,78,24,28.44,5521,0,Miranda,1,1,Fiber Optic,40.210895,-123.86,0,53.5,0,0,Offer B,867,1,0,0,0,57,0,0.0,1621.0800000000004,0.0,3035.8,0,1,95553
2980,0,0,0,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.45,1866.45,0,39,0,6.75,4118,0,Myers Flat,0,0,NA,40.267158,-123.80591299999999,0,25.45,0,0,Offer A,644,0,0,0,0,72,0,0.0,486.0,0.0,1866.45,0,0,95554
2981,1,0,0,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.5,1430.95,0,24,0,47.31,4416,0,Orick,0,1,NA,41.336354,-124.044354,0,20.5,0,0,Offer A,494,0,0,0,0,67,1,0.0,3169.77,0.0,1430.95,1,0,95555
2982,1,0,1,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.85,1071.6,0,47,0,39.48,4886,0,Orleans,0,1,NA,41.269521000000005,-123.546958,1,20.85,3,2,Offer B,574,0,0,1,0,52,0,0.0,2052.96,0.0,1071.6,0,0,95556
2983,1,0,1,1,71,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.9,6457.15,0,57,27,31.33,4444,0,Petrolia,1,1,Fiber Optic,40.274302,-124.210902,1,89.9,3,6,Offer A,300,1,0,1,1,71,0,1743.0,2224.43,0.0,6457.15,0,0,95558
2984,0,0,1,0,26,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,26.0,684.05,0,56,0,33.47,2244,0,Phillipsville,0,0,NA,40.184094,-123.74548700000001,1,26.0,0,7,None,163,0,1,1,0,26,1,0.0,870.22,0.0,684.05,0,0,95559
2985,0,0,0,0,35,1,1,Fiber optic,1,1,1,1,Two year,1,Mailed check,113.2,3914.05,0,49,8,30.5,5723,0,Redway,1,0,Fiber Optic,40.142256,-123.85292700000001,0,113.2,0,0,None,1851,1,0,0,1,35,0,0.0,1067.5,0.0,3914.05,0,1,95560
2986,0,0,1,1,55,1,0,Fiber optic,0,0,0,0,Two year,1,Credit card (automatic),69.05,3842.6,0,52,17,27.87,4318,0,Rio Dell,0,0,Fiber Optic,40.485849,-124.163234,1,69.05,2,3,Offer B,3284,0,0,1,0,55,1,653.0,1532.85,0.0,3842.6,0,0,95562
2987,0,0,1,1,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.1,670.35,0,61,0,24.27,3700,0,Salyer,0,0,NA,40.89866,-123.539754,1,20.1,3,2,None,660,0,1,1,0,33,1,0.0,800.91,0.0,670.35,0,0,95563
2988,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,109.65,7880.25,0,20,73,6.89,6181,0,Samoa,1,1,DSL,40.809636,-124.189977,1,109.65,0,2,Offer A,395,0,0,1,1,72,1,0.0,496.08,0.0,7880.25,1,1,95564
2989,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.2,19.2,0,37,0,17.89,3383,0,Scotia,0,1,NA,40.440636,-124.098739,0,19.2,3,0,None,1125,0,0,0,0,1,0,0.0,17.89,0.0,19.2,0,0,95565
2990,1,0,0,0,10,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Mailed check,33.9,298.45,1,42,33,0.0,2529,1,Smith River,0,1,DSL,41.950683000000005,-124.097094,0,35.256,0,0,None,2020,0,0,0,1,10,2,98.0,0.0,0.0,298.45,0,0,95567
2991,0,1,1,0,37,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,90.0,3371.75,0,66,19,15.6,4048,0,Somes Bar,1,0,Fiber Optic,41.444606,-123.47189499999999,1,90.0,0,8,None,202,1,2,1,0,37,1,641.0,577.1999999999998,0.0,3371.75,0,0,95568
2992,1,0,0,0,12,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Mailed check,34.0,442.45,0,35,6,0.0,3215,0,Redcrest,0,1,DSL,40.363446,-123.83504099999999,0,34.0,0,0,Offer D,400,1,0,0,0,12,0,0.0,0.0,0.0,442.45,0,1,95569
2993,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.4,20.4,0,27,0,27.5,4540,0,Trinidad,0,1,NA,41.162295,-124.027381,1,20.4,2,3,None,2369,0,0,1,0,1,3,0.0,27.5,0.0,20.4,1,0,95570
2994,1,0,1,0,62,0,No phone service,DSL,1,1,0,0,Two year,1,Credit card (automatic),38.6,2345.55,0,56,29,0.0,4558,0,Weott,0,1,Fiber Optic,40.310119,-123.909449,1,38.6,0,8,Offer B,270,1,0,1,0,62,2,680.0,0.0,0.0,2345.55,0,0,95571
2995,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),25.25,25.25,0,40,15,0.0,4831,0,Willow Creek,0,0,DSL,40.949011999999996,-123.655847,0,25.25,0,0,Offer E,1666,0,0,0,0,1,2,0.0,0.0,0.0,25.25,0,1,95573
2996,0,0,0,0,18,1,1,DSL,1,0,0,0,Month-to-month,1,Mailed check,60.6,1156.35,0,64,9,10.97,4459,0,Leggett,1,0,Fiber Optic,39.873371,-123.741474,0,60.6,0,0,Offer D,321,0,0,0,0,18,0,0.0,197.46,0.0,1156.35,0,1,95585
2997,1,1,1,0,69,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.95,6143.15,1,65,4,16.34,6363,1,Piercy,0,1,Cable,39.955587,-123.681175,1,93.54799999999999,0,1,None,200,0,1,1,0,69,6,0.0,1127.46,6.79,6143.15,0,1,95587
2998,1,0,0,0,2,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.75,144.8,0,19,52,43.56,4545,0,Fallbrook,0,1,DSL,33.362575,-117.299644,0,74.75,0,0,Offer E,42239,0,0,0,0,2,0,75.0,87.12,0.0,144.8,1,0,92028
2999,1,0,1,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.6,414.95,0,43,0,4.7,2276,0,Zenia,0,1,NA,40.170357,-123.417298,1,20.6,2,6,Offer D,259,0,1,1,0,19,3,0.0,89.3,0.0,414.95,0,0,95595
3000,1,0,0,0,12,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.45,1059.55,1,41,25,12.36,3330,1,Amador City,0,1,Fiber Optic,38.431407,-120.8421,0,87.82799999999999,0,0,None,222,0,0,0,0,12,4,265.0,148.32,0.0,1059.55,0,0,95601
3001,1,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,181.8,0,36,0,13.72,5380,0,Auburn,0,1,NA,38.99003,-121.11440800000001,0,20.4,0,0,Offer E,18197,0,0,0,0,9,0,0.0,123.48,0.0,181.8,0,0,95602
3002,1,0,0,0,27,1,0,DSL,1,0,1,1,One year,0,Electronic check,81.7,2212.55,0,58,4,49.25,2445,0,Auburn,1,1,Fiber Optic,38.912881,-121.08276599999999,0,81.7,0,0,None,24944,1,0,0,1,27,1,89.0,1329.75,0.0,2212.55,0,0,95603
3003,1,0,0,1,27,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,79.5,2180.55,1,35,32,24.72,2518,1,West Sacramento,0,1,Cable,38.592745,-121.54003600000001,0,82.68,0,0,None,12756,1,0,0,0,27,2,698.0,667.4399999999998,0.0,2180.55,0,0,95605
3004,1,0,1,1,1,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Mailed check,89.15,89.15,1,44,20,32.35,3123,1,Brooks,0,1,Cable,38.809804,-122.24138300000001,1,92.716,0,1,None,382,0,3,1,1,1,3,0.0,32.35,0.0,89.15,0,1,95606
3005,0,1,0,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.3,459.95,0,78,0,18.39,3740,0,Capay,0,0,NA,38.681651,-122.130569,0,20.3,0,0,None,262,0,0,0,0,24,2,0.0,441.36,0.0,459.95,0,0,95607
3006,1,1,0,0,14,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.95,1036.75,1,67,12,16.32,2075,1,Carmichael,0,1,Cable,38.626128,-121.328011,0,77.94800000000002,0,0,Offer D,58830,0,0,0,0,14,2,124.0,228.48,39.29,1036.75,0,0,95608
3007,0,1,0,0,32,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.4,2276.95,1,70,10,33.22,2091,1,Citrus Heights,0,0,Cable,38.69508,-121.271616,0,77.376,0,0,Offer C,43718,0,1,0,0,32,3,228.0,1063.04,44.31,2276.95,0,0,95610
3008,0,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.0,211.95,0,31,0,46.49,3731,0,Clarksburg,0,0,NA,38.384648,-121.578701,0,20.0,0,0,Offer D,1417,0,1,0,0,11,1,0.0,511.39,0.0,211.95,0,0,95612
3009,1,0,0,0,1,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,25.0,25,0,41,0,3.39,2371,0,Cool,0,1,NA,38.880621999999995,-120.97386499999999,0,25.0,0,0,Offer E,3674,0,0,0,0,1,0,0.0,3.39,0.0,25.0,0,0,95614
3010,1,1,0,1,38,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,80.45,3162.65,0,76,27,45.13,2926,0,Courtland,0,1,Fiber Optic,38.311609000000004,-121.554034,0,80.45,2,0,None,699,0,0,0,0,38,0,85.39,1714.94,0.0,3162.65,0,1,95615
3011,0,0,1,1,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,210.65,0,45,0,16.13,2427,0,Davis,0,0,NA,38.508734999999994,-121.67881299999999,1,19.75,2,6,Offer E,67411,0,0,1,0,9,1,0.0,145.17,0.0,210.65,0,0,95616
3012,1,0,1,1,54,1,1,DSL,1,1,0,0,Two year,1,Credit card (automatic),65.65,3566.7,0,25,52,24.59,5725,0,Davis,0,1,DSL,38.544002,-121.68555900000001,1,65.65,2,1,Offer B,648,1,0,1,0,54,2,1855.0,1327.86,0.0,3566.7,1,0,95618
3013,0,0,0,0,29,1,1,DSL,0,0,1,1,One year,1,Credit card (automatic),71.0,2080.1,0,47,4,41.38,4226,0,Diamond Springs,0,0,Cable,38.683605,-120.811852,0,71.0,0,0,None,4426,0,0,0,1,29,0,83.0,1200.02,0.0,2080.1,0,0,95619
3014,1,1,1,0,44,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,89.2,4040.2,0,72,30,14.65,2925,0,Dixon,1,1,Fiber Optic,38.392821000000005,-121.799917,1,89.2,0,6,Offer B,18529,0,0,1,0,44,0,1212.0,644.6,0.0,4040.2,0,0,95620
3015,1,0,1,1,59,1,0,DSL,1,1,1,1,Two year,1,Electronic check,86.75,5186,0,21,73,42.37,5020,0,Citrus Heights,1,1,Fiber Optic,38.69549,-121.307864,1,86.75,3,4,Offer B,41636,1,0,1,1,59,2,3786.0,2499.83,0.0,5186.0,1,0,95621
3016,0,0,0,0,3,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.3,196.15,1,45,8,25.96,3190,1,El Dorado,0,0,Fiber Optic,38.63153,-120.84260900000001,0,57.512,0,0,None,4097,0,1,0,1,3,4,16.0,77.88,0.0,196.15,0,0,95623
3017,0,0,1,1,18,1,0,DSL,1,1,0,0,One year,1,Mailed check,61.5,1087.45,0,22,51,40.36,3479,0,Elk Grove,0,0,Fiber Optic,38.434138,-121.30587,1,61.5,2,7,Offer D,38534,1,0,1,0,18,2,555.0,726.48,0.0,1087.45,1,0,95624
3018,1,1,0,0,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.1,1672.15,0,73,0,14.69,6388,0,Elmira,0,1,NA,38.349195,-121.902943,0,25.1,0,0,None,171,0,1,0,0,67,3,0.0,984.23,0.0,1672.15,0,0,95625
3019,0,0,1,1,22,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,55.15,1206.05,1,32,21,5.26,5115,1,Elverta,0,0,Cable,38.734997,-121.463719,1,57.356,1,1,None,6197,1,0,1,0,22,0,0.0,115.72,0.0,1206.05,0,1,95626
3020,1,0,0,1,33,0,No phone service,DSL,1,0,0,0,One year,0,Credit card (automatic),34.05,1113.95,0,64,12,0.0,3044,0,Esparto,0,1,Fiber Optic,38.834469,-122.12719299999999,0,34.05,2,0,None,2756,1,0,0,0,33,1,0.0,0.0,0.0,1113.95,0,1,95627
3021,1,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,107.05,0,31,0,24.16,4281,0,Fair Oaks,0,1,NA,38.652065,-121.25441000000001,0,19.95,0,0,None,40750,0,0,0,0,5,0,0.0,120.8,0.0,107.05,0,0,95628
3022,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,38.15,0,33,0,34.57,4079,0,Fiddletown,0,0,NA,38.513484000000005,-120.704613,0,19.95,0,0,Offer E,850,0,0,0,0,2,0,0.0,69.14,0.0,38.15,0,0,95629
3023,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.7,6339.3,0,25,30,33.75,4193,0,Folsom,1,1,Cable,38.672638,-121.147403,1,89.7,1,10,Offer A,51855,1,0,1,1,72,0,0.0,2430.0,0.0,6339.3,1,1,95630
3024,1,0,0,1,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,184.1,0,34,0,45.83,4195,0,Foresthill,0,1,NA,39.031876000000004,-120.81114099999999,0,20.4,2,0,Offer E,5714,0,0,0,0,9,0,0.0,412.47,0.0,184.1,0,0,95631
3025,1,0,1,1,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,26.3,1688.9,0,54,0,14.54,6066,0,Galt,0,1,NA,38.274451,-121.259201,1,26.3,2,2,Offer A,24194,0,0,1,0,67,1,0.0,974.18,0.0,1688.9,0,0,95632
3026,0,0,1,0,16,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.95,1378.25,1,34,8,6.82,3075,1,Garden Valley,0,0,DSL,38.852544,-120.83766899999999,1,88.348,0,1,None,2536,0,1,1,0,16,5,0.0,109.12,0.0,1378.25,0,1,95633
3027,0,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.7,137.6,0,59,0,26.47,3330,0,Georgetown,0,0,NA,38.9386,-120.78551399999999,0,20.7,0,0,Offer E,2723,0,0,0,0,8,1,0.0,211.76,0.0,137.6,0,0,95634
3028,1,0,0,0,5,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Mailed check,43.25,219,1,30,65,0.0,5824,1,Greenwood,1,1,Fiber Optic,38.921333000000004,-120.897718,0,44.98,0,0,None,1140,1,3,0,0,5,4,0.0,0.0,0.0,219.0,0,1,95635
3029,1,0,1,1,23,1,1,DSL,0,0,0,0,One year,1,Credit card (automatic),48.35,1067.15,1,60,13,5.8,4580,1,Grizzly Flats,0,1,Fiber Optic,38.636102,-120.522149,1,50.284000000000006,0,1,None,659,0,0,1,0,23,0,139.0,133.4,0.0,1067.15,0,0,95636
3030,1,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.55,79.55,1,59,7,4.04,5593,1,Guinda,0,1,DSL,38.830739,-122.196202,0,82.73200000000001,0,0,None,228,0,0,0,0,1,4,0.0,4.04,0.0,79.55,0,0,95637
3031,0,1,1,0,50,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.05,3444.85,1,69,26,4.6,5746,1,Herald,0,0,DSL,38.313447,-121.12388600000001,1,73.892,0,1,None,1745,0,0,1,0,50,5,896.0,230.0,0.0,3444.85,0,0,95638
3032,1,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.45,369.05,0,50,0,39.34,5347,0,Hood,0,1,NA,38.375325,-121.507935,0,19.45,0,0,Offer D,213,0,0,0,0,17,1,0.0,668.7800000000002,0.0,369.05,0,0,95639
3033,0,0,1,0,68,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),110.8,7553.6,0,61,14,46.7,4545,0,Ione,1,0,Fiber Optic,38.33788,-120.954202,1,110.8,0,2,Offer A,9752,0,0,1,1,68,3,0.0,3175.600000000001,0.0,7553.6,0,1,95640
3034,1,0,0,0,1,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,84.5,84.5,1,31,13,6.89,4340,1,Isleton,0,1,Fiber Optic,38.154823,-121.601358,0,87.88000000000002,0,0,None,2010,0,0,0,0,1,3,0.0,6.89,0.0,84.5,0,0,95641
3035,0,1,1,0,25,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.3,1813.1,0,75,24,38.59,4442,0,Jackson,0,0,Fiber Optic,38.336216,-120.76901000000001,1,69.3,0,7,None,6202,0,0,1,0,25,0,0.0,964.75,0.0,1813.1,0,1,95642
3036,1,0,0,0,67,0,No phone service,DSL,1,0,1,0,One year,1,Bank transfer (automatic),49.35,3321.35,0,30,85,0.0,5905,0,Knights Landing,1,1,DSL,38.875508,-121.76586599999999,0,49.35,0,0,Offer A,1793,1,0,0,0,67,1,0.0,0.0,0.0,3321.35,0,1,95645
3037,1,0,0,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.35,707.5,0,20,0,36.78,2433,0,Kirkwood,0,1,NA,38.631489,-120.01516699999999,0,20.35,0,0,None,129,0,0,0,0,32,3,0.0,1176.96,0.0,707.5,1,0,95646
3038,0,1,1,0,67,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,105.6,7112.15,0,74,10,11.91,5768,0,Lincoln,0,0,Fiber Optic,38.922812,-121.312005,1,105.6,0,3,None,15286,0,0,1,1,67,0,711.0,797.97,0.0,7112.15,0,0,95648
3039,1,1,1,0,72,0,No phone service,DSL,1,1,1,1,Two year,1,Credit card (automatic),64.45,4641.1,0,76,9,0.0,5295,0,Loomis,1,1,Cable,38.809175,-121.171375,1,64.45,0,9,None,11191,1,0,1,1,72,0,0.0,0.0,0.0,4641.1,0,1,95650
3040,1,0,1,0,71,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),108.6,7690.9,1,57,12,5.76,4982,1,Lotus,1,1,Fiber Optic,38.815515000000005,-120.916997,1,112.944,0,1,Offer A,485,1,2,1,1,71,2,923.0,408.96,0.0,7690.9,0,0,95651
3041,1,0,0,1,1,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,49.9,49.9,0,29,76,6.35,3239,0,Madison,0,1,DSL,38.674276,-121.96186599999999,0,49.9,1,0,Offer E,844,0,0,0,0,1,0,0.0,6.35,0.0,49.9,1,1,95653
3042,1,0,0,0,46,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),30.3,1380.1,1,57,29,0.0,2243,1,Mather,0,1,DSL,38.549822,-121.266725,0,31.511999999999997,0,0,None,929,0,4,0,0,46,3,400.0,0.0,0.0,1380.1,0,0,95655
3043,0,1,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,30.4,78.65,1,73,14,0.0,4002,1,Newcastle,1,0,DSL,38.883224,-121.15918,0,31.616,0,0,None,6096,0,0,0,0,2,3,11.0,0.0,0.0,78.65,0,0,95658
3044,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.4,45.4,1,32,29,38.31,2168,1,Nicolaus,0,0,Fiber Optic,38.788897999999996,-121.608624,0,47.216,0,0,None,751,0,4,0,0,1,1,0.0,38.31,0.0,45.4,0,0,95659
3045,0,0,1,0,48,1,0,DSL,0,1,0,1,One year,1,Electronic check,65.65,3094.65,0,27,42,49.88,5427,0,North Highlands,1,0,DSL,38.671295,-121.388251,1,65.65,0,6,Offer B,32202,0,1,1,1,48,2,0.0,2394.24,0.0,3094.65,1,1,95660
3046,0,0,1,0,61,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),103.3,6518.35,0,63,22,18.03,5401,0,Roseville,1,0,DSL,38.736684999999994,-121.25198400000001,1,103.3,0,6,Offer B,25173,1,0,1,1,61,2,143.4,1099.8300000000004,0.0,6518.35,0,1,95661
3047,0,0,1,0,32,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Bank transfer (automatic),84.15,2585.95,1,53,14,37.48,4017,1,Orangevale,0,0,Cable,38.689174,-121.21843500000001,1,87.516,0,1,None,32040,0,1,1,1,32,3,362.0,1199.36,0.0,2585.95,0,0,95662
3048,0,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.45,82.7,0,22,59,18.7,5694,0,Penryn,0,0,DSL,38.859093,-121.182872,0,44.45,0,0,Offer E,2048,0,0,0,0,2,1,49.0,37.4,0.0,82.7,1,0,95663
3049,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.75,58.85,1,41,0,24.63,2647,1,Pilot Hill,0,0,NA,38.803731,-121.04379899999999,0,19.75,0,0,Offer E,1173,0,0,0,0,3,2,0.0,73.89,0.0,58.85,0,0,95664
3050,0,0,0,0,5,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),85.4,425.9,1,62,19,43.51,3716,1,Pine Grove,0,0,Fiber Optic,38.400264,-120.641274,0,88.816,0,0,Offer E,4354,1,0,0,1,5,6,81.0,217.55,0.0,425.9,0,0,95665
3051,0,0,1,1,71,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),89.9,6342.7,0,22,85,37.57,5835,0,Pioneer,1,0,DSL,38.546999,-120.27111399999998,1,89.9,1,9,Offer A,5501,1,0,1,1,71,0,0.0,2667.47,0.0,6342.7,1,1,95666
3052,1,0,1,0,37,1,1,DSL,1,0,0,0,Month-to-month,1,Mailed check,55.05,2030.75,0,57,10,27.41,3839,0,Placerville,0,1,Fiber Optic,38.733714,-120.79521299999999,1,55.05,0,6,None,34146,0,0,1,0,37,0,0.0,1014.17,0.0,2030.75,0,1,95667
3053,1,0,1,1,65,1,1,Fiber optic,0,0,1,1,Two year,1,Bank transfer (automatic),104.1,6700.05,0,40,57,39.52,4024,0,Pleasant Grove,1,1,Fiber Optic,38.833554,-121.498102,1,104.1,3,0,Offer B,901,1,0,0,1,65,1,0.0,2568.8,0.0,6700.05,0,1,95668
3054,0,0,0,1,67,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),106.6,7244.7,0,19,59,18.74,5895,0,Plymouth,0,0,Cable,38.489273,-120.89161399999999,0,106.6,2,0,Offer A,2220,1,0,0,1,67,0,0.0,1255.58,0.0,7244.7,1,1,95669
3055,1,0,0,1,49,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),75.2,3678.3,1,62,26,19.08,5283,1,Rancho Cordova,0,1,Cable,38.602723,-121.279913,0,78.20800000000001,0,0,None,49729,0,0,0,0,49,3,956.0,934.92,0.0,3678.3,0,0,95670
3056,1,0,1,1,50,1,1,DSL,1,0,1,0,Two year,1,Credit card (automatic),70.5,3486.65,0,53,28,44.49,4022,0,Rescue,0,1,Fiber Optic,38.724321999999994,-120.99123700000001,1,70.5,2,10,Offer B,3815,1,0,1,0,50,0,0.0,2224.5,0.0,3486.65,0,1,95672
3057,1,0,1,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.6,411.15,0,43,0,15.76,2888,0,Rio Linda,0,1,NA,38.688764,-121.457596,1,19.6,2,1,None,14010,0,0,1,0,25,1,0.0,394.0,0.0,411.15,0,0,95673
3058,0,0,0,1,17,1,1,DSL,0,0,0,0,One year,1,Mailed check,55.85,937.5,1,50,23,24.31,5472,1,Rio Oso,1,0,Cable,38.954144,-121.48253600000001,0,58.083999999999996,0,0,None,947,0,0,0,0,17,0,0.0,413.27,0.0,937.5,0,1,95674
3059,0,0,1,1,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.05,1559.15,0,45,0,17.93,4582,0,River Pines,0,0,NA,38.545775,-120.743325,1,24.05,3,5,Offer B,364,0,0,1,0,64,0,0.0,1147.52,0.0,1559.15,0,0,95675
3060,1,0,1,0,25,0,No phone service,DSL,0,0,1,0,One year,1,Credit card (automatic),38.1,970.4,0,37,24,0.0,2315,0,Rocklin,1,1,Fiber Optic,38.7904,-121.23697299999999,1,38.1,0,10,None,21510,0,0,1,0,25,0,0.0,0.0,0.0,970.4,0,1,95677
3061,1,1,0,0,23,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.4,2483.5,1,74,32,17.62,5507,1,Roseville,1,1,Cable,38.759751,-121.288545,0,110.656,0,0,None,30614,0,0,0,0,23,0,795.0,405.2600000000001,0.0,2483.5,0,0,95678
3062,1,1,1,0,24,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,34.25,828.2,0,68,28,0.0,2525,0,Sheridan,1,1,DSL,38.984756,-121.345074,1,34.25,0,3,None,1219,1,0,1,0,24,0,0.0,0.0,0.0,828.2,0,1,95681
3063,0,0,0,0,37,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.05,3810.55,0,64,22,17.46,2904,0,Shingle Springs,1,0,DSL,38.598936,-120.96309199999999,0,100.05,0,0,Offer C,24738,0,0,0,1,37,1,838.0,646.02,0.0,3810.55,0,0,95682
3064,0,0,0,0,21,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,68.65,1493.2,0,60,11,30.59,2006,0,Sloughhouse,0,0,DSL,38.470423,-121.114897,0,68.65,0,0,Offer D,4731,0,0,0,0,21,2,164.0,642.39,0.0,1493.2,0,0,95683
3065,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.8,45.8,0,34,21,13.62,2614,0,Somerset,0,1,DSL,38.606703,-120.58665900000001,0,45.8,0,0,None,2958,0,0,0,0,1,0,0.0,13.62,0.0,45.8,0,1,95684
3066,0,0,0,0,10,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,75.75,777.3,0,37,21,39.85,4525,0,Sutter Creek,0,0,Cable,38.432145,-120.77068999999999,0,75.75,0,0,None,4610,0,0,0,0,10,4,163.0,398.5,0.0,777.3,0,0,95685
3067,1,0,0,0,6,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,84.4,556.35,1,53,10,21.97,4539,1,Thornton,0,1,Fiber Optic,38.157794,-121.520223,0,87.77600000000002,0,0,None,1472,0,2,0,1,6,2,56.0,131.82,0.0,556.35,0,0,95686
3068,1,0,1,0,51,1,1,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),96.4,4911.05,0,63,8,35.0,4745,0,Vacaville,0,1,Fiber Optic,38.333133000000004,-121.920151,1,96.4,0,7,Offer B,63157,0,0,1,1,51,1,0.0,1785.0,0.0,4911.05,0,1,95687
3069,0,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.55,187.35,0,63,0,4.76,3595,0,Vacaville,0,0,NA,38.419088,-122.02456799999999,0,20.55,0,0,None,32564,0,0,0,0,10,1,0.0,47.6,0.0,187.35,0,0,95688
3070,0,0,0,0,6,0,No phone service,DSL,1,1,0,1,Month-to-month,0,Credit card (automatic),50.95,307.6,0,43,23,0.0,3474,0,Volcano,0,0,Fiber Optic,38.481902000000005,-120.603668,0,50.95,0,0,Offer E,1273,1,0,0,1,6,1,0.0,0.0,0.0,307.6,0,1,95689
3071,1,0,1,1,47,1,1,DSL,1,1,1,1,Two year,1,Mailed check,90.5,4318.35,0,30,48,11.74,3413,0,Walnut Grove,1,1,DSL,38.240419,-121.587535,1,90.5,3,10,Offer B,2344,1,0,1,1,47,1,0.0,551.78,0.0,4318.35,0,1,95690
3072,0,0,1,1,61,1,1,DSL,1,1,0,1,One year,1,Electronic check,79.4,4820.55,0,52,20,40.48,4666,0,West Sacramento,1,0,Cable,38.627951,-121.59328700000002,1,79.4,2,3,Offer B,19050,1,0,1,1,61,0,0.0,2469.28,0.0,4820.55,0,1,95691
3073,0,0,0,0,52,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),58.75,3038.55,0,40,19,0.0,5122,0,Wheatland,1,0,Cable,39.043387,-121.40983700000001,0,58.75,0,0,Offer B,3600,0,0,0,1,52,2,0.0,0.0,0.0,3038.55,0,1,95692
3074,0,0,1,1,35,1,1,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),59.45,2136.9,0,42,23,39.11,3682,0,Wilton,0,0,Fiber Optic,38.392559000000006,-121.22509299999999,1,59.45,3,0,Offer C,5889,0,0,0,0,35,2,49.15,1368.85,0.0,2136.9,0,1,95693
3075,1,0,1,0,71,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),105.7,7472.15,0,52,28,29.11,4420,0,Winters,1,1,DSL,38.578604,-122.024579,1,105.7,0,8,Offer A,8406,0,0,1,1,71,0,0.0,2066.81,0.0,7472.15,0,1,95694
3076,0,0,0,0,6,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,56.25,389.1,1,44,24,17.18,4110,1,Woodland,0,0,Cable,38.71967,-121.862416,0,58.5,0,0,Offer E,38547,0,0,0,0,6,4,0.0,103.08,0.0,389.1,0,1,95695
3077,1,0,1,0,45,1,0,DSL,1,0,0,0,Two year,0,Credit card (automatic),53.3,2296.25,0,37,4,43.27,2929,0,Alta,1,1,DSL,39.218096,-120.79153000000001,1,53.3,0,10,None,751,0,1,1,0,45,3,0.0,1947.15,0.0,2296.25,0,1,95701
3078,0,1,0,0,2,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.55,187.45,1,78,28,5.49,5512,1,Applegate,0,0,Cable,38.983388,-120.98881399999999,0,88.97200000000001,0,0,Offer E,1526,0,0,0,0,2,0,52.0,10.98,0.0,187.45,0,0,95703
3079,0,0,0,0,4,1,0,DSL,0,1,1,1,Month-to-month,1,Bank transfer (automatic),68.65,261.25,1,51,25,10.64,5274,1,Camino,0,0,DSL,38.748315999999996,-120.67551200000001,0,71.39600000000002,0,0,Offer E,4829,0,0,0,1,4,6,65.0,42.56,0.0,261.25,0,0,95709
3080,1,0,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,24.3,38.45,0,19,59,0.0,2515,0,Colfax,0,1,Cable,39.084645,-120.89401399999998,0,24.3,0,0,Offer E,8525,0,0,0,0,2,2,23.0,0.0,0.0,38.45,1,0,95713
3081,1,0,0,0,4,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,77.85,299.2,1,48,31,42.8,2140,1,Dutch Flat,0,1,Cable,39.197215,-120.83679,0,80.964,0,0,Offer E,350,0,0,0,0,4,2,93.0,171.2,0.0,299.2,0,0,95714
3082,1,0,0,0,51,1,1,DSL,1,0,0,0,One year,0,Credit card (automatic),59.9,3043.6,0,59,3,9.85,5233,0,Emigrant Gap,0,1,Fiber Optic,39.23754,-120.720196,0,59.9,0,0,None,185,1,0,0,0,51,0,91.0,502.35,0.0,3043.6,0,0,95715
3083,1,0,1,1,60,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),23.95,1506.4,0,37,0,28.45,5449,0,Gold Run,0,1,NA,39.170376,-120.838404,1,23.95,2,1,None,407,0,0,1,0,60,1,0.0,1707.0,0.0,1506.4,0,0,95717
3084,1,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.15,163.7,0,40,0,48.61,4004,0,Kyburz,0,1,NA,38.766036,-120.209673,0,20.15,0,0,Offer E,183,0,0,0,0,9,1,0.0,437.49,0.0,163.7,0,0,95720
3085,1,0,0,0,3,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),105.35,323.25,1,50,15,13.83,3662,1,Echo Lake,1,1,Cable,38.851842,-120.076204,0,109.564,0,0,Offer E,69,0,0,0,1,3,3,0.0,41.49,0.0,323.25,0,1,95721
3086,1,0,0,0,17,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),95.65,1640,0,58,5,21.14,3139,0,Meadow Vista,1,1,DSL,39.003358,-121.022539,0,95.65,0,0,None,3747,1,0,0,1,17,0,82.0,359.38,0.0,1640.0,0,0,95722
3087,0,0,0,0,8,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,87.05,762.1,1,48,9,45.59,2545,1,Pollock Pines,0,0,Cable,38.733908,-120.45341599999999,0,90.53200000000001,0,0,Offer E,8577,0,1,0,0,8,3,69.0,364.72,0.0,762.1,0,0,95726
3088,1,0,1,1,46,1,0,DSL,1,0,1,1,Two year,0,Mailed check,81.0,3846.35,0,37,10,45.95,4280,0,Soda Springs,1,1,Cable,39.279068,-120.414275,1,81.0,1,1,None,88,1,0,1,1,46,3,0.0,2113.7000000000007,0.0,3846.35,0,1,95728
3089,0,0,0,0,68,1,0,DSL,1,1,1,1,Two year,1,Credit card (automatic),82.45,5646.6,0,21,59,14.86,5308,0,Twin Bridges,1,0,DSL,38.805481,-120.13287,0,82.45,0,0,Offer A,25,1,1,0,1,68,1,0.0,1010.48,0.0,5646.6,1,1,95735
3090,1,0,0,0,1,1,0,DSL,0,0,1,0,Month-to-month,1,Mailed check,53.5,53.5,1,22,80,14.58,5094,1,Weimar,0,1,Fiber Optic,39.00978,-120.978273,0,55.64,0,0,None,31,0,0,0,0,1,0,0.0,14.58,0.0,53.5,1,0,95736
3091,0,0,1,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.5,79.05,0,52,0,44.73,3233,0,Rancho Cordova,0,0,NA,38.591134000000004,-121.161585,1,20.5,0,8,None,299,0,0,1,0,4,1,0.0,178.92,0.0,79.05,0,0,95742
3092,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,25.1,25.1,1,35,31,0.0,4769,1,Granite Bay,0,0,Cable,38.749466,-121.184196,0,26.104000000000006,0,0,None,20675,0,1,0,0,1,5,0.0,0.0,0.0,25.1,0,1,95746
3093,1,0,0,1,28,1,0,DSL,0,1,0,0,One year,1,Credit card (automatic),54.4,1516.6,0,55,22,34.43,4711,0,Roseville,0,1,Fiber Optic,38.784329,-121.373245,0,54.4,1,0,Offer C,25418,1,0,0,0,28,1,334.0,964.04,0.0,1516.6,0,0,95747
3094,0,0,0,0,39,1,0,DSL,0,1,1,0,One year,1,Credit card (automatic),58.6,2224.5,0,23,58,48.17,5662,0,Elk Grove,0,0,Fiber Optic,38.353629999999995,-121.44195,0,58.6,0,0,Offer C,47065,0,0,0,0,39,1,0.0,1878.63,0.0,2224.5,1,1,95758
3095,1,0,0,0,11,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,84.8,888.75,0,54,15,30.57,4924,0,El Dorado Hills,1,1,Fiber Optic,38.684437,-121.05563400000001,0,84.8,0,0,None,22028,0,0,0,1,11,1,133.0,336.27,0.0,888.75,0,0,95762
3096,0,0,1,0,71,0,No phone service,DSL,0,1,1,1,Two year,1,Credit card (automatic),61.4,4310.35,0,46,27,0.0,5119,0,Rocklin,1,0,Cable,38.823278,-121.281856,1,61.4,0,2,Offer A,15494,1,0,1,1,71,0,0.0,0.0,0.0,4310.35,0,1,95765
3097,1,0,0,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,42.9,0,42,0,49.53,3000,0,Woodland,0,1,NA,38.694081,-121.69443100000001,0,20.4,2,0,None,15022,0,0,0,0,2,0,0.0,99.06,0.0,42.9,0,0,95776
3098,1,1,1,0,30,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,79.65,2365.15,1,77,4,6.23,2174,1,Sacramento,1,1,Cable,38.584505,-121.491956,1,82.83600000000001,0,1,Offer C,16599,0,0,1,0,30,5,95.0,186.9,0.0,2365.15,0,0,95814
3099,0,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.15,353.65,0,35,0,4.38,4650,0,Sacramento,0,0,NA,38.608405,-121.449942,0,20.15,0,0,None,25355,0,0,0,0,17,0,0.0,74.46,0.0,353.65,0,0,95815
3100,0,0,1,0,55,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),94.45,5073.1,0,64,16,34.61,5577,0,Sacramento,1,0,Fiber Optic,38.574856,-121.46503999999999,1,94.45,0,1,None,16164,0,0,1,0,55,1,812.0,1903.55,0.0,5073.1,0,0,95816
3101,0,0,0,0,58,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),79.8,4526.85,0,47,14,22.71,5709,0,Sacramento,0,0,Cable,38.550722,-121.457314,0,79.8,0,0,None,14966,0,0,0,0,58,1,0.0,1317.18,0.0,4526.85,0,1,95817
3102,0,0,0,0,5,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,54.2,308.25,1,21,76,3.61,5476,1,Sacramento,0,0,Cable,38.556306,-121.49581699999999,0,56.368,0,0,None,21313,1,0,0,0,5,0,0.0,18.05,0.0,308.25,1,1,95818
3103,0,1,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.45,19.45,1,70,0,22.92,3848,1,Sacramento,0,0,NA,38.567594,-121.43750700000001,0,19.45,0,0,None,15975,0,0,0,0,1,1,0.0,22.92,0.0,19.45,0,0,95819
3104,1,1,0,0,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.05,678.45,0,66,25,39.77,2003,0,Sacramento,0,1,Fiber Optic,38.53508,-121.444144,0,74.05,0,0,Offer E,37031,0,0,0,0,9,3,170.0,357.93,0.0,678.45,0,0,95820
3105,1,0,0,0,26,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),49.15,1237.3,0,36,8,44.11,2752,0,Sacramento,0,1,DSL,38.625096,-121.38365800000001,0,49.15,0,0,Offer C,35426,1,0,0,0,26,3,0.0,1146.86,0.0,1237.3,0,1,95821
3106,0,0,0,0,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.4,1023.95,0,36,0,12.62,6233,0,Sacramento,0,0,NA,38.512569,-121.49518400000001,0,19.4,0,0,None,44683,0,0,0,0,50,2,0.0,631.0,0.0,1023.95,0,0,95822
3107,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),113.65,8182.75,0,35,22,29.0,5411,0,Sacramento,1,0,DSL,38.475465,-121.443625,1,113.65,0,10,Offer A,72199,1,2,1,1,72,1,1800.0,2088.0,0.0,8182.75,0,0,95823
3108,0,0,0,1,43,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),106.0,4532.3,0,47,10,10.19,3528,0,Sacramento,0,0,DSL,38.517295000000004,-121.439819,0,106.0,2,0,None,30580,1,0,0,1,43,0,0.0,438.17,0.0,4532.3,0,1,95824
3109,1,0,0,0,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.95,1444.05,0,52,0,47.82,4246,0,Sacramento,0,1,NA,38.590035,-121.41245500000001,0,25.95,0,0,None,30715,0,0,0,0,56,0,0.0,2677.92,0.0,1444.05,0,0,95825
3110,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.1,19.1,0,28,0,5.02,3313,0,Sacramento,0,0,NA,38.542532,-121.378826,0,19.1,0,0,None,38818,0,0,0,0,1,0,0.0,5.02,0.0,19.1,1,0,95826
3111,1,0,1,1,72,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,103.4,7372.65,1,47,25,3.07,5055,1,Sacramento,1,1,Cable,38.549184999999994,-121.32838600000001,1,107.53600000000002,0,1,None,19611,0,0,1,1,72,2,1843.0,221.04,0.0,7372.65,0,0,95827
3112,1,0,1,0,72,1,1,Fiber optic,1,1,0,1,Two year,1,Bank transfer (automatic),100.55,7325.1,0,62,15,43.84,6082,0,Sacramento,0,1,Fiber Optic,38.486938,-121.39580500000001,1,100.55,0,5,Offer A,54880,1,0,1,1,72,1,1099.0,3156.4800000000005,0.0,7325.1,0,0,95828
3113,1,0,1,0,36,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.4,3474.2,0,58,12,40.58,5111,0,Sacramento,0,1,Fiber Optic,38.486502,-121.334051,1,95.4,0,4,Offer C,11396,0,0,1,1,36,0,0.0,1460.88,0.0,3474.2,0,1,95829
3114,1,0,0,0,5,1,0,DSL,0,0,1,1,Month-to-month,0,Bank transfer (automatic),75.15,392.65,0,51,4,45.69,5900,0,Sacramento,1,1,DSL,38.490508,-121.284171,0,75.15,0,0,None,592,1,0,0,1,5,1,0.0,228.45,0.0,392.65,0,1,95830
3115,0,0,0,0,13,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,84.45,1058.6,1,60,4,21.88,5801,1,Sacramento,1,0,DSL,38.494832,-121.52944699999999,0,87.82799999999999,0,0,None,42832,0,0,0,0,13,2,42.0,284.44,0.0,1058.6,0,0,95831
3116,0,1,0,0,44,1,0,Fiber optic,0,1,0,1,One year,0,Credit card (automatic),89.15,3990.75,0,70,19,35.39,4368,0,Sacramento,1,0,DSL,38.445939,-121.49685500000001,0,89.15,0,0,Offer B,9063,0,2,0,1,44,1,758.0,1557.16,0.0,3990.75,0,0,95832
3117,0,1,1,1,70,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,107.9,7475.85,0,65,17,9.4,5899,0,Sacramento,1,0,Fiber Optic,38.619049,-121.517552,1,107.9,2,2,None,31422,1,1,1,1,70,2,1271.0,658.0,0.0,7475.85,0,0,95833
3118,1,0,0,0,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.5,835.5,0,60,0,18.14,4220,0,Sacramento,0,1,NA,38.646209000000006,-121.52446,0,19.5,0,0,None,8403,0,0,0,0,44,1,0.0,798.1600000000002,0.0,835.5,0,0,95834
3119,0,1,1,0,32,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),85.95,2628.6,1,78,10,48.95,2431,1,Sacramento,0,0,Cable,38.685069,-121.543709,1,89.38799999999999,0,0,Offer C,854,0,0,0,0,32,7,263.0,1566.4,0.0,2628.6,0,0,95835
3120,0,0,1,0,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.95,1718.35,0,23,0,45.12,4106,0,Sacramento,0,0,NA,38.691607,-121.60228400000001,1,24.95,0,10,None,264,0,0,1,0,69,0,0.0,3113.28,0.0,1718.35,1,0,95837
3121,0,1,0,0,16,1,0,DSL,0,0,1,0,Month-to-month,0,Electronic check,59.4,1023.9,1,75,18,36.83,5556,1,Sacramento,0,0,DSL,38.646096,-121.44243300000001,0,61.776,0,0,None,34894,1,1,0,0,16,3,0.0,589.28,0.0,1023.9,0,1,95838
3122,1,1,1,1,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.5,1193.55,0,73,0,35.14,5443,0,Sacramento,0,1,NA,38.660441999999996,-121.346321,1,19.5,1,8,None,20993,0,0,1,0,68,2,0.0,2389.52,0.0,1193.55,0,0,95841
3123,1,0,0,0,16,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),69.95,1205.5,0,43,27,27.43,5596,0,Sacramento,0,1,Fiber Optic,38.687367,-121.34848000000001,0,69.95,0,0,None,31373,0,0,0,0,16,1,0.0,438.88,0.0,1205.5,0,1,95842
3124,1,0,1,1,68,1,0,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),82.85,5776.45,0,52,27,27.59,5184,0,Antelope,0,1,Cable,38.715498,-121.36341100000001,1,82.85,1,1,None,36432,1,0,1,1,68,0,0.0,1876.12,0.0,5776.45,0,1,95843
3125,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.0,78.9,0,31,0,20.16,3022,0,Sacramento,0,1,NA,38.585826000000004,-121.376263,0,19.0,0,0,None,23362,0,0,0,0,4,1,0.0,80.64,0.0,78.9,0,0,95864
3126,0,0,1,1,26,0,No phone service,DSL,1,1,0,0,Month-to-month,0,Credit card (automatic),38.85,1025.15,0,40,23,0.0,3970,0,Marysville,0,0,Fiber Optic,39.19514,-121.503883,1,38.85,3,4,Offer C,38091,1,0,1,0,26,0,236.0,0.0,0.0,1025.15,0,0,95901
3127,0,0,0,0,29,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,30.6,856.35,1,53,8,0.0,3615,1,Beale Afb,0,0,Cable,39.125310999999996,-121.392283,0,31.824,0,0,None,5654,0,3,0,0,29,5,69.0,0.0,0.0,856.35,0,0,95903
3128,1,0,0,1,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.35,122,0,39,0,8.01,3161,0,Alleghany,0,1,NA,39.467828000000004,-120.84138600000001,0,20.35,1,0,None,118,0,1,0,0,5,4,0.0,40.05,0.0,122.0,0,0,95910
3129,1,0,1,0,70,1,1,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),95.0,6602.9,0,48,16,31.13,6259,0,Arbuckle,1,1,Cable,38.982372999999995,-122.047751,1,95.0,0,5,None,4796,0,0,1,0,70,0,1056.0,2179.1,0.0,6602.9,0,0,95912
3130,1,0,1,0,24,1,0,DSL,1,0,1,1,One year,0,Bank transfer (automatic),74.4,1712.9,0,61,30,32.86,4310,0,Bangor,0,1,Fiber Optic,39.396584999999995,-121.38028999999999,1,74.4,0,10,Offer C,626,1,0,1,1,24,2,0.0,788.64,0.0,1712.9,0,1,95914
3131,0,1,1,0,72,1,1,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),78.45,5682.25,0,68,13,15.82,4032,0,Berry Creek,1,0,Fiber Optic,39.657228,-121.37778,1,78.45,0,10,None,1279,1,0,1,1,72,1,0.0,1139.04,0.0,5682.25,0,1,95916
3132,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.3,74.3,0,37,21,39.55,3063,0,Biggs,0,1,Cable,39.457388,-121.818201,0,74.3,0,0,None,3169,1,0,0,0,1,0,0.0,39.55,0.0,74.3,0,1,95917
3133,1,0,1,0,70,0,No phone service,DSL,0,1,0,1,One year,1,Bank transfer (automatic),51.05,3635.15,0,19,41,0.0,4042,0,Browns Valley,1,1,Fiber Optic,39.292334000000004,-121.32059699999999,1,51.05,0,10,None,1477,1,0,1,1,70,0,1490.0,0.0,0.0,3635.15,1,0,95918
3134,0,0,1,1,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.2,702.9,0,56,0,20.57,3043,0,Brownsville,0,0,NA,39.440687,-121.26358300000001,1,19.2,2,3,Offer C,1237,0,0,1,0,36,3,0.0,740.52,0.0,702.9,0,0,95919
3135,0,1,0,0,38,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.55,3734.25,1,75,2,47.39,3474,1,Butte City,0,0,Cable,39.449794,-121.93637199999999,0,103.53200000000001,0,0,Offer C,303,1,1,0,0,38,2,0.0,1800.82,0.0,3734.25,0,1,95920
3136,0,0,0,0,17,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.0,1144.5,1,51,19,7.66,4390,1,Camptonville,0,0,Fiber Optic,39.432127,-121.09928700000002,0,72.8,0,0,None,632,0,1,0,0,17,2,217.0,130.22,0.0,1144.5,0,0,95922
3137,0,0,1,1,41,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),109.1,4454.25,0,28,59,20.41,4854,0,Canyon Dam,1,0,Fiber Optic,40.171312,-121.120605,1,109.1,2,3,None,86,1,0,1,1,41,1,2628.0,836.8100000000002,0.0,4454.25,1,0,95923
3138,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.3,45.3,1,37,29,26.41,2293,1,Challenge,0,0,Cable,39.461768,-121.195825,0,47.111999999999995,0,0,None,262,0,1,0,0,1,1,0.0,26.41,0.0,45.3,0,0,95925
3139,1,0,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),29.85,75.6,1,64,12,0.0,4268,1,Chico,0,1,Fiber Optic,39.745712,-121.84333000000001,0,31.044000000000004,0,0,None,35808,1,0,0,0,2,0,9.0,0.0,0.0,75.6,0,0,95926
3140,1,0,0,0,14,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,76.45,1117.55,0,20,26,18.46,2292,0,Chico,1,1,Cable,39.681488,-121.83721000000001,0,76.45,0,0,None,32848,0,0,0,0,14,0,0.0,258.44,0.0,1117.55,1,1,95928
3141,1,1,0,0,2,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),95.1,180.25,1,76,22,12.96,4486,1,Clipper Mills,1,1,Cable,39.562239,-121.14836000000001,0,98.904,0,0,Offer E,282,1,0,0,0,2,4,0.0,25.92,0.0,180.25,0,1,95930
3142,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.8,19.8,1,40,0,9.66,5600,1,Colusa,0,1,NA,39.273096,-122.05076299999999,0,19.8,0,0,None,7503,0,0,0,0,1,4,0.0,9.66,0.0,19.8,0,0,95932
3143,1,0,1,1,13,1,1,DSL,0,1,1,0,Month-to-month,1,Electronic check,72.8,930.05,0,33,23,13.77,2862,0,Crescent Mills,1,1,Fiber Optic,40.080342,-120.95780500000001,1,72.8,2,4,None,178,1,0,1,0,13,1,21.39,179.01,0.0,930.05,0,1,95934
3144,1,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,18.95,110.15,0,24,0,27.54,5920,0,Dobbins,0,1,NA,39.381174,-121.21191,0,18.95,0,0,None,614,0,0,0,0,6,2,0.0,165.24,0.0,110.15,1,0,95935
3145,0,0,0,0,4,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),76.65,333.6,1,36,19,24.09,4580,1,Downieville,0,0,Cable,39.578792,-120.780786,0,79.71600000000002,0,0,None,404,0,0,0,0,4,3,63.0,96.36,0.0,333.6,0,0,95936
3146,0,0,1,1,5,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Mailed check,99.15,465.05,1,45,28,9.23,2283,1,Dunnigan,0,0,Cable,38.931425,-121.946081,1,103.116,0,1,None,19,1,0,1,1,5,2,130.0,46.15000000000001,0.0,465.05,0,0,95937
3147,0,0,1,0,15,1,0,Fiber optic,1,0,1,1,Month-to-month,0,Electronic check,101.75,1669.4,0,55,13,24.12,2919,0,Durham,1,0,Cable,39.607831,-121.77795900000001,1,101.75,0,8,None,3524,0,0,1,1,15,2,217.0,361.8,0.0,1669.4,0,0,95938
3148,0,0,0,0,47,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Credit card (automatic),75.45,3545.1,0,19,69,48.03,4995,0,Elk Creek,0,0,Fiber Optic,39.53222,-122.594879,0,75.45,0,0,None,587,0,0,0,0,47,0,244.61,2257.41,0.0,3545.1,1,1,95939
3149,0,0,0,0,8,1,0,DSL,0,0,0,1,Month-to-month,0,Mailed check,64.1,504.05,0,19,73,45.04,2804,0,Forbestown,1,0,Fiber Optic,39.531028000000006,-121.24807,0,64.1,0,0,None,452,1,0,0,1,8,0,368.0,360.32,0.0,504.05,1,0,95941
3150,1,0,0,0,17,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,25.65,440.2,0,63,11,0.0,3090,0,Forest Ranch,0,1,DSL,40.077028000000006,-121.49416799999999,0,25.65,0,0,None,1351,0,0,0,0,17,0,48.0,0.0,0.0,440.2,0,0,95942
3151,1,0,1,1,15,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Mailed check,75.1,1151.55,0,39,17,32.73,4634,0,Glenn,0,1,DSL,39.597975,-122.032248,1,75.1,1,7,None,1454,0,0,1,0,15,2,0.0,490.94999999999993,0.0,1151.55,0,1,95943
3152,0,0,0,0,26,1,0,Fiber optic,1,0,0,1,One year,1,Bank transfer (automatic),95.85,2475.35,0,60,4,40.14,3834,0,Goodyears Bar,1,0,Fiber Optic,39.564113,-120.86883600000002,0,95.85,0,0,Offer C,76,1,0,0,1,26,2,0.0,1043.64,0.0,2475.35,0,1,95944
3153,0,0,0,0,23,1,1,DSL,1,0,0,0,Month-to-month,0,Electronic check,54.4,1249.25,0,40,11,48.63,2989,0,Grass Valley,0,0,Fiber Optic,39.194539,-120.98806599999999,0,54.4,0,0,None,23990,0,0,0,0,23,1,0.0,1118.49,0.0,1249.25,0,1,95945
3154,0,1,0,0,4,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,72.75,317.75,0,76,8,35.67,4503,0,Penn Valley,0,0,Cable,39.203817,-121.19583999999999,0,72.75,0,0,None,9752,0,0,0,0,4,0,25.0,142.68,0.0,317.75,0,0,95946
3155,1,0,0,1,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.85,535.05,0,54,0,2.0,2941,0,Greenville,0,1,NA,40.160385999999995,-120.83542800000001,0,19.85,3,0,Offer C,2064,0,0,0,0,29,1,0.0,58.0,0.0,535.05,0,0,95947
3156,0,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.05,461.3,0,50,0,30.28,2692,0,Gridley,0,0,NA,39.346897999999996,-121.75953700000001,0,19.05,0,0,Offer C,9763,0,0,0,0,25,0,0.0,757.0,0.0,461.3,0,0,95948
3157,1,0,0,0,9,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.95,431,1,57,29,2.88,5023,1,Grass Valley,0,1,Fiber Optic,39.099204,-121.13796200000002,0,46.74800000000001,0,0,Offer E,17922,0,2,0,0,9,4,125.0,25.92,0.0,431.0,0,0,95949
3158,1,0,1,0,18,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,49.55,878.35,1,53,29,19.05,2815,1,Grimes,1,1,DSL,39.033058000000004,-121.89571799999999,1,51.532,0,1,None,531,0,1,1,0,18,5,0.0,342.9000000000001,0.0,878.35,0,1,95950
3159,1,1,0,0,3,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.85,335.75,0,65,28,37.78,4496,0,Hamilton City,0,1,Cable,39.732766999999996,-122.042298,0,94.85,0,0,Offer E,1931,0,2,0,1,3,1,0.0,113.34,0.0,335.75,0,1,95951
3160,0,0,1,1,69,0,No phone service,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),46.25,3121.4,0,29,69,0.0,4180,0,Live Oak,1,0,Fiber Optic,39.258746,-121.77696999999999,1,46.25,2,10,None,8695,1,0,1,0,69,0,215.38,0.0,0.0,3121.4,1,1,95953
3161,1,0,0,0,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.35,324.8,0,24,0,26.02,2400,0,Magalia,0,1,NA,39.933852,-121.58437099999999,0,19.35,0,0,Offer D,11168,0,0,0,0,14,0,0.0,364.28,0.0,324.8,1,0,95954
3162,1,0,0,0,19,1,1,DSL,0,0,1,1,Month-to-month,0,Mailed check,69.6,1394.55,0,54,4,13.76,3349,0,Maxwell,0,1,Cable,39.281194,-122.226568,0,69.6,0,0,Offer D,1146,0,0,0,1,19,0,0.0,261.44,0.0,1394.55,0,1,95955
3163,1,1,0,0,39,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,90.7,3413.25,0,76,3,20.06,5028,0,Meadow Valley,0,1,DSL,39.937017,-121.058043,0,90.7,0,0,None,301,0,0,0,1,39,0,0.0,782.3399999999998,0.0,3413.25,0,1,95956
3164,1,0,0,0,31,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.4,3143.65,0,20,76,19.38,2025,0,Meridian,1,1,Cable,39.068071,-121.83263799999999,0,101.4,0,0,Offer C,776,0,0,0,1,31,2,2389.0,600.78,0.0,3143.65,1,0,95957
3165,1,0,1,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.25,439.75,0,61,0,40.81,3000,0,Nevada City,0,1,NA,39.333737,-120.858667,1,20.25,2,5,Offer C,17269,0,0,1,0,24,0,0.0,979.44,0.0,439.75,0,0,95959
3166,1,0,1,0,14,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),48.8,664.4,0,39,24,21.34,2168,0,North San Juan,0,1,DSL,39.423046,-120.984472,1,48.8,0,4,Offer D,565,1,0,1,0,14,0,159.0,298.76,0.0,664.4,0,0,95960
3167,0,0,1,0,64,1,0,DSL,1,1,0,1,Two year,1,Mailed check,74.35,4759.55,0,23,42,18.03,4781,0,Olivehurst,1,0,Fiber Optic,39.082568,-121.55325,1,74.35,0,2,None,6439,1,0,1,1,64,1,0.0,1153.92,0.0,4759.55,1,1,95961
3168,0,0,0,0,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.35,1033,0,29,0,17.88,5247,0,Oregon House,0,0,NA,39.342587,-121.24983300000001,0,19.35,0,0,None,1519,0,0,0,0,50,0,0.0,894.0,29.5,1033.0,1,0,95962
3169,1,0,1,1,52,1,0,DSL,0,1,1,0,One year,1,Electronic check,68.75,3482.85,0,45,19,5.51,4172,0,Orland,1,1,Fiber Optic,39.748037,-122.30216899999999,1,68.75,2,9,None,13706,1,0,1,0,52,0,662.0,286.52,16.86,3482.85,0,0,95963
3170,1,0,0,0,28,1,1,Fiber optic,0,1,1,1,One year,0,Electronic check,100.2,2688.45,0,31,13,12.36,5137,0,Oroville,0,1,DSL,39.624561,-121.552866,0,100.2,0,0,Offer C,17782,0,1,0,1,28,3,0.0,346.08,42.64,2688.45,0,1,95965
3171,0,0,0,0,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.85,435.25,0,40,0,22.29,5422,0,Oroville,0,0,NA,39.473896,-121.415927,0,20.85,0,0,Offer D,28382,0,0,0,0,21,0,0.0,468.09,1.31,435.25,0,0,95966
3172,1,0,0,1,25,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,95.9,2448.75,1,55,4,5.27,2241,1,Palermo,0,1,Cable,39.435756,-121.552071,0,99.736,0,0,None,1254,0,0,0,1,25,1,0.0,131.75,0.0,2448.75,0,1,95968
3173,0,0,1,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.35,307,0,33,0,1.64,2185,0,Paradise,0,0,NA,39.69676,-121.644379,1,19.35,0,3,Offer D,28318,0,0,1,0,17,2,0.0,27.88,10.57,307.0,0,0,95969
3174,1,0,1,0,58,0,No phone service,DSL,0,0,1,1,One year,1,Credit card (automatic),45.0,2689.35,0,53,23,0.0,5006,0,Princeton,0,1,Fiber Optic,39.424957,-122.03930700000001,1,45.0,0,0,None,495,0,0,0,1,58,3,0.0,0.0,0.0,2689.35,0,1,95970
3175,1,1,1,0,17,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Bank transfer (automatic),81.5,1329.2,1,70,18,9.5,3443,1,Quincy,0,1,Fiber Optic,39.971228,-121.04116599999999,1,84.76,0,1,None,6189,0,2,1,0,17,1,239.0,161.5,0.0,1329.2,0,0,95971
3176,0,0,1,0,51,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.5,1281.25,0,59,0,20.47,5447,0,Chico,0,0,NA,39.903271999999994,-121.843567,1,25.5,0,7,None,26971,0,0,1,0,51,0,0.0,1043.97,0.0,1281.25,0,0,95973
3177,1,0,1,1,72,0,No phone service,DSL,1,0,1,0,Two year,0,Mailed check,48.9,3527,0,53,53,0.0,5415,0,Richvale,1,1,Cable,39.495768,-121.747472,1,48.9,3,3,None,74,1,0,1,0,72,0,1869.0,0.0,34.44,3527.0,0,0,95974
3178,1,0,1,0,52,1,0,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,84.1,4348.65,1,40,15,38.37,6216,1,Rough And Ready,0,1,Fiber Optic,39.225634,-121.15616299999999,1,87.464,0,1,None,1601,0,0,1,0,52,0,652.0,1995.24,0.0,4348.65,0,0,95975
3179,0,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.6,561.15,0,62,0,15.41,2896,0,Smartville,0,0,NA,39.176595,-121.291692,0,19.6,0,0,None,963,0,1,0,0,27,1,0.0,416.07,13.07,561.15,0,0,95977
3180,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,63.6,0,38,0,40.2,4258,0,Stirling City,0,0,NA,39.904002,-121.527823,0,20.0,0,0,None,28,0,0,0,0,3,0,0.0,120.6,0.0,63.6,0,0,95978
3181,0,0,1,0,64,1,1,DSL,1,1,0,1,Two year,1,Mailed check,81.3,5129.3,0,33,4,16.61,5254,0,Stonyford,1,0,DSL,39.288127,-122.41584099999999,1,81.3,0,6,None,844,1,0,1,1,64,0,0.0,1063.04,22.34,5129.3,0,1,95979
3182,0,0,1,0,45,1,0,Fiber optic,0,0,1,1,Two year,1,Credit card (automatic),95.2,4285.8,0,51,18,48.02,3363,0,Strawberry Valley,0,0,Fiber Optic,39.584579999999995,-121.09325600000001,1,95.2,0,3,None,101,1,0,1,1,45,1,0.0,2160.9,43.95,4285.8,0,1,95981
3183,1,1,1,0,3,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Mailed check,36.45,93.7,1,67,22,0.0,3766,1,Sutter,0,1,Cable,39.172777,-121.80584499999999,1,37.908,0,1,Offer E,3193,0,3,1,0,3,1,21.0,0.0,0.0,93.7,0,0,95982
3184,0,0,1,0,71,1,1,DSL,0,1,1,1,Two year,1,Credit card (automatic),83.3,5894.5,0,56,18,13.41,4264,0,Taylorsville,1,0,Fiber Optic,40.053684000000004,-120.74311599999999,1,83.3,0,9,None,513,1,1,1,1,71,3,0.0,952.11,37.44,5894.5,0,1,95983
3185,0,1,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,25.05,25.05,1,69,23,0.0,4842,1,Twain,0,0,DSL,40.022184,-121.06238400000001,0,26.052000000000003,0,0,Offer E,73,0,2,0,0,1,4,0.0,0.0,0.0,25.05,0,1,95984
3186,0,0,1,1,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.3,1160.75,0,35,0,17.21,4424,0,Washington,0,0,NA,39.34128,-120.78686699999999,1,20.3,1,6,None,145,0,0,1,0,58,1,0.0,998.18,25.57,1160.75,0,0,95986
3187,1,0,1,1,34,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.85,3091.75,0,25,85,18.36,3096,0,Williams,1,1,Fiber Optic,39.117537,-122.284654,1,89.85,3,5,None,4579,0,0,1,0,34,0,2628.0,624.24,14.93,3091.75,1,0,95987
3188,0,0,0,0,8,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.85,365.55,1,48,28,37.79,2269,1,Willows,0,0,Fiber Optic,39.493990999999994,-122.286363,0,51.843999999999994,0,0,None,8812,0,0,0,0,8,4,0.0,302.32,13.01,365.55,0,1,95988
3189,0,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.8,272.95,0,49,0,17.43,4167,0,Yuba City,0,0,NA,39.027409999999996,-121.61498200000001,1,19.8,1,4,Offer D,34967,0,0,1,0,15,2,0.0,261.45,18.55,272.95,0,0,95991
3190,1,0,1,1,66,0,No phone service,DSL,0,0,1,1,Two year,0,Bank transfer (automatic),54.65,3632,0,49,28,0.0,4051,0,Yuba City,1,1,Cable,39.075694,-121.70606000000001,1,54.65,3,0,None,27786,1,0,0,1,66,0,1017.0,0.0,46.75,3632.0,0,0,95993
3191,1,1,0,0,12,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),29.35,381.2,0,79,4,0.0,3606,0,Redding,0,1,Fiber Optic,40.587919,-122.46473200000001,0,29.35,0,0,None,31586,0,0,0,0,12,0,0.0,0.0,38.98,381.2,0,1,96001
3192,1,0,0,0,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.15,1035.5,0,49,0,29.31,6339,0,Redding,0,1,NA,40.527834000000006,-122.318749,0,19.15,0,0,None,30338,0,0,0,0,58,0,0.0,1699.98,28.7,1035.5,0,0,96002
3193,0,0,1,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.1,52,0,32,0,45.33,3863,0,Redding,0,0,NA,40.677649,-122.29467,1,19.1,2,9,None,41476,0,0,1,0,3,1,0.0,135.99,0.0,52.0,0,0,96003
3194,0,1,1,0,43,0,No phone service,DSL,0,1,1,1,Month-to-month,0,Credit card (automatic),55.55,2342.2,1,70,23,0.0,2573,1,Adin,1,0,Fiber Optic,41.171578000000004,-120.91316100000002,1,57.772,0,1,Offer B,615,0,1,1,0,43,2,0.0,0.0,0.0,2342.2,0,1,96006
3195,0,0,0,0,9,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,80.55,653.9,0,38,13,32.57,3581,0,Anderson,1,0,DSL,40.448632,-122.306657,0,80.55,0,0,None,21418,0,0,0,0,9,1,8.5,293.13,2.28,653.9,0,1,96007
3196,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.25,71.2,0,60,0,1.47,4331,0,Bella Vista,0,0,NA,40.722733000000005,-122.10966599999999,0,20.25,0,0,None,899,0,0,0,0,3,0,0.0,4.41,0.0,71.2,0,0,96008
3197,0,0,1,1,22,1,0,DSL,0,1,1,1,One year,1,Bank transfer (automatic),69.5,1498.2,1,22,84,35.04,5922,1,Bieber,0,0,Fiber Optic,41.083464,-121.107929,1,72.28,0,1,None,595,0,0,1,1,22,3,125.85,770.88,49.57,1498.2,1,1,96009
3198,1,0,1,0,40,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),106.0,4178.65,0,37,28,29.46,5118,0,Big Bar,1,1,Fiber Optic,40.775271999999994,-123.28741399999998,1,106.0,0,1,Offer B,269,0,0,1,1,40,0,0.0,1178.4,47.02,4178.65,0,1,96010
3199,0,0,0,0,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.5,1821.8,0,50,0,9.82,5182,0,Big Bend,0,0,NA,41.096569,-121.87908200000001,0,25.5,0,0,None,265,0,1,0,0,68,2,0.0,667.76,16.85,1821.8,0,0,96011
3200,1,0,1,0,54,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.3,5278.15,1,47,25,35.46,4019,1,Burney,1,1,Cable,40.946785,-121.719489,1,108.47200000000001,0,1,None,4552,0,1,1,1,54,2,0.0,1914.84,11.45,5278.15,0,1,96013
3201,0,0,0,0,50,1,1,DSL,0,1,1,1,Two year,1,Mailed check,79.6,4024.2,0,39,14,48.45,5592,0,Callahan,0,0,DSL,41.388397,-122.79463600000001,0,79.6,0,0,Offer B,290,1,0,0,1,50,0,563.0,2422.5,0.0,4024.2,0,0,96014
3202,1,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.25,55.25,0,21,69,39.19,3255,0,Canby,0,1,DSL,41.486953,-120.913975,0,55.25,0,0,None,417,0,0,0,1,1,1,0.0,39.19,0.0,55.25,1,1,96015
3203,0,0,1,0,72,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),88.05,6520.8,0,49,24,38.28,6247,0,Cassel,1,0,Cable,40.936285,-121.57269199999999,1,88.05,0,1,None,344,1,0,1,1,72,0,156.5,2756.16,29.11,6520.8,0,1,96016
3204,1,0,0,1,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.4,854.9,0,58,0,26.41,3200,0,Castella,0,1,NA,41.121108,-122.33661299999999,0,20.4,3,0,Offer B,228,0,0,0,0,40,1,0.0,1056.4,32.55,854.9,0,0,96017
3205,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),117.6,8308.9,0,28,48,47.02,6173,0,Shasta Lake,1,0,Fiber Optic,40.692523,-122.369876,1,117.6,1,10,None,6277,1,0,1,1,72,2,0.0,3385.44,5.44,8308.9,1,1,96019
3206,0,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,109.2,0,60,0,47.46,3142,0,Chester,0,0,NA,40.243494,-121.15473300000001,0,20.0,0,0,None,2664,0,0,0,0,6,1,0.0,284.76,0.0,109.2,0,0,96020
3207,0,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.65,92.05,0,62,0,41.93,2878,0,Corning,0,0,NA,39.913777,-122.289984,0,19.65,0,0,None,13840,0,0,0,0,5,2,0.0,209.65,0.0,92.05,0,0,96021
3208,1,0,1,0,48,1,1,DSL,0,1,0,1,One year,1,Credit card (automatic),70.55,3420.5,0,41,8,38.82,3997,0,Cottonwood,1,1,Cable,40.336392,-122.44853300000001,1,70.55,0,7,Offer B,12348,0,2,1,1,48,1,274.0,1863.36,0.0,3420.5,0,0,96022
3209,0,0,0,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.85,93.85,1,49,13,16.15,3014,1,Dorris,0,0,Fiber Optic,41.949216,-122.05006200000001,0,97.604,0,0,Offer E,1162,0,0,0,1,1,1,0.0,16.15,0.0,93.85,0,1,96023
3210,0,0,1,1,64,1,0,DSL,1,0,1,0,One year,0,Mailed check,65.8,4068,0,39,17,26.7,4754,0,Douglas City,0,0,Fiber Optic,40.586588,-122.903677,1,65.8,2,5,Offer B,960,1,0,1,0,64,1,692.0,1708.8,27.79,4068.0,0,0,96024
3211,0,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.05,337.9,0,63,0,3.84,4828,0,Dunsmuir,0,0,NA,41.212695000000004,-122.392067,0,20.05,0,0,Offer D,2602,0,0,0,0,17,1,0.0,65.28,43.68,337.9,0,0,96025
3212,1,0,1,0,40,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.0,3168.75,0,41,27,39.22,2478,0,Etna,1,1,Fiber Optic,41.405193,-123.008567,1,80.0,0,8,Offer B,2156,0,0,1,0,40,1,0.0,1568.8,41.74,3168.75,0,1,96027
3213,0,0,1,1,41,0,No phone service,DSL,1,0,0,0,One year,0,Credit card (automatic),35.4,1412.4,0,37,16,0.0,4375,0,Fall River Mills,1,0,Fiber Optic,41.017282,-121.46894499999999,1,35.4,2,1,Offer B,1902,0,0,1,0,41,0,0.0,0.0,0.0,1412.4,0,1,96028
3214,1,1,0,0,51,1,1,Fiber optic,0,1,0,0,One year,1,Bank transfer (automatic),79.6,3974.7,0,69,11,24.92,4673,0,Flournoy,0,1,DSL,39.847840000000005,-122.544556,0,79.6,0,0,None,84,0,0,0,0,51,2,0.0,1270.92,16.73,3974.7,0,1,96029
3215,1,0,1,0,41,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.25,3439,0,36,3,39.39,5757,0,Forks Of Salmon,0,1,DSL,41.232128,-123.194748,1,80.25,0,10,Offer B,170,0,0,1,0,41,2,103.0,1614.99,2.18,3439.0,0,0,96031
3216,0,0,1,1,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.45,50.45,1,47,32,9.73,2426,1,Escondido,1,0,Cable,33.141265000000004,-116.967221,1,52.468,2,1,Offer E,48690,0,0,1,0,1,2,0.0,9.73,0.0,50.45,0,1,92027
3217,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.45,42.45,0,31,0,47.19,2606,0,French Gulch,0,0,NA,40.740138,-122.587476,0,20.45,0,0,None,373,0,0,0,0,2,3,0.0,94.38,0.0,42.45,0,0,96033
3218,1,0,0,0,68,1,0,Fiber optic,0,1,0,0,One year,0,Credit card (automatic),79.6,5461.45,0,50,21,18.53,5210,0,Gazelle,1,1,DSL,41.411315,-122.697236,0,79.6,0,0,None,392,0,0,0,0,68,1,1147.0,1260.04,3.26,5461.45,0,0,96034
3219,0,0,1,1,24,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.7,571.75,0,42,0,20.74,5302,0,Gerber,0,0,NA,40.031940000000006,-122.176023,1,24.7,3,7,None,3357,0,0,1,0,24,0,0.0,497.76,0.0,571.75,0,0,96035
3220,1,0,1,0,70,1,1,DSL,1,0,0,1,Two year,0,Credit card (automatic),77.3,5498.2,0,22,41,4.8,6252,0,Greenview,1,1,Fiber Optic,41.528541,-122.955018,1,77.3,0,2,None,295,1,0,1,1,70,0,2254.0,336.0,26.87,5498.2,1,0,96037
3221,1,0,0,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,29.75,96.85,0,58,18,0.0,3425,0,Grenada,0,1,Cable,41.599978,-122.539381,0,29.75,0,0,Offer E,616,1,0,0,0,3,1,17.0,0.0,0.0,96.85,0,0,96038
3222,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),44.9,111.05,0,56,17,5.08,4370,0,Happy Camp,0,1,Fiber Optic,41.831901,-123.487478,0,44.9,0,0,None,1294,0,0,0,0,2,1,0.0,10.16,0.0,111.05,0,1,96039
3223,1,0,1,0,3,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Credit card (automatic),29.8,94.4,0,62,4,0.0,5614,0,Hat Creek,0,1,DSL,40.789799,-121.474529,1,29.8,0,1,Offer E,397,0,0,1,0,3,1,4.0,0.0,0.0,94.4,0,0,96040
3224,0,0,0,0,7,1,1,DSL,0,0,1,1,Month-to-month,1,Electronic check,74.65,521.1,1,33,21,48.82,4612,1,Fallbrook,0,0,Fiber Optic,33.362575,-117.299644,0,77.63600000000002,0,0,Offer E,42239,1,0,0,1,7,1,109.0,341.74,28.35,521.1,0,0,92028
3225,0,0,0,0,13,1,0,DSL,1,0,1,1,Month-to-month,1,Electronic check,71.95,923.85,0,54,5,10.66,3605,0,Hornbrook,0,0,Fiber Optic,41.962127,-122.52769599999999,0,71.95,0,0,Offer D,1026,0,0,0,1,13,2,46.0,138.58,10.47,923.85,0,0,96044
3226,1,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.75,141.1,0,44,0,47.19,4476,0,Hyampom,0,1,NA,40.648024,-123.465088,0,20.75,0,0,Offer E,268,0,1,0,0,7,1,0.0,330.33,0.0,141.1,0,0,96046
3227,1,0,1,1,12,1,0,DSL,0,0,1,0,Month-to-month,1,Mailed check,56.3,628.65,0,49,29,17.27,2047,0,Igo,0,1,Fiber Optic,40.524535,-122.647172,1,56.3,2,5,Offer D,911,0,0,1,0,12,0,0.0,207.24,0.0,628.65,0,1,96047
3228,1,0,1,1,53,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,105.25,5576.3,0,40,27,3.78,6365,0,Junction City,1,1,Fiber Optic,40.913191999999995,-123.06597,1,105.25,1,7,Offer B,734,0,1,1,1,53,3,1506.0,200.34,0.0,5576.3,0,0,96048
3229,0,0,0,0,12,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.2,1046.1,1,53,26,12.75,3975,1,Klamath River,0,0,Cable,41.816595,-122.94828700000001,0,97.96799999999999,0,0,None,482,0,0,0,1,12,4,272.0,153.0,7.39,1046.1,0,0,96050
3230,1,0,1,1,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.55,1245.6,0,48,0,10.67,6002,0,Lakehead,0,1,NA,40.883853,-122.41825800000001,1,19.55,2,4,Offer B,1236,0,1,1,0,63,2,0.0,672.21,0.0,1245.6,0,0,96051
3231,0,0,0,0,15,1,0,DSL,1,1,1,1,Month-to-month,0,Mailed check,84.45,1287.85,0,58,2,8.97,4653,0,Lewiston,1,0,DSL,40.704293,-122.803899,0,84.45,0,0,Offer D,1845,1,0,0,1,15,0,26.0,134.55,0.0,1287.85,0,0,96052
3232,1,0,1,1,36,1,0,DSL,1,1,0,0,One year,0,Mailed check,53.65,1939.35,0,40,19,8.0,4113,0,Lookout,0,1,DSL,41.280478,-121.160249,1,53.65,1,2,None,386,0,0,1,0,36,0,0.0,288.0,0.0,1939.35,0,1,96054
3233,1,1,1,0,4,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,29.9,118.25,0,78,5,0.0,2914,0,Los Molinos,1,1,Cable,40.059385,-122.091481,1,29.9,0,3,Offer E,3756,0,1,1,0,4,1,0.59,0.0,0.0,118.25,0,1,96055
3234,0,0,1,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.7,452.55,0,51,0,30.41,4642,0,Mcarthur,0,0,NA,41.108309999999996,-121.36036200000001,1,19.7,1,8,None,1554,0,0,1,0,24,1,0.0,729.84,0.0,452.55,0,0,96056
3235,0,0,0,0,61,0,No phone service,DSL,1,1,0,0,One year,0,Credit card (automatic),43.7,2696.55,0,59,8,0.0,4051,0,Mccloud,1,0,DSL,41.251321999999995,-122.105209,0,43.7,0,0,Offer B,1586,1,0,0,0,61,0,216.0,0.0,0.0,2696.55,0,0,96057
3236,1,0,0,0,16,1,1,DSL,0,1,0,0,Month-to-month,0,Electronic check,55.3,875.35,0,43,4,5.79,3771,0,Macdoel,0,1,DSL,41.769709000000006,-121.92063,0,55.3,0,0,None,816,0,0,0,0,16,2,35.0,92.64,0.0,875.35,0,0,96058
3237,1,0,1,1,65,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.85,1267.05,0,55,0,33.47,6009,0,Manton,0,1,NA,40.426679,-121.850421,1,19.85,1,5,Offer B,598,0,0,1,0,65,2,0.0,2175.55,0.0,1267.05,0,0,96059
3238,0,0,1,1,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.65,494.9,0,40,0,12.71,4184,0,Mill Creek,0,0,NA,40.331975,-121.460674,1,19.65,2,4,None,78,0,0,1,0,26,0,0.0,330.4600000000001,0.0,494.9,0,0,96061
3239,1,0,0,0,16,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,49.45,799,0,29,59,48.45,3446,0,Millville,0,1,Cable,40.531257000000004,-122.14813899999999,0,49.45,0,0,None,830,1,0,0,0,16,0,0.0,775.2,0.0,799.0,1,1,96062
3240,0,0,1,0,54,1,1,Fiber optic,1,1,1,1,One year,0,Bank transfer (automatic),106.55,5763.3,1,59,23,8.83,4893,1,Mineral,0,0,Cable,40.408796,-121.579609,1,110.81200000000001,0,2,None,124,0,0,1,1,54,0,132.56,476.82,0.0,5763.3,0,1,96063
3241,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.1,20.1,1,33,0,16.81,5747,1,Fallbrook,0,1,NA,33.362575,-117.299644,0,20.1,0,0,Offer E,42239,0,0,0,0,1,0,0.0,16.81,0.0,20.1,0,0,92028
3242,1,0,0,1,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.45,106.9,0,19,0,29.15,3353,0,Montgomery Creek,0,1,NA,40.877552,-121.885884,0,20.45,1,0,Offer E,431,0,0,0,0,5,0,0.0,145.75,0.0,106.9,1,0,96065
3243,0,0,0,0,19,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Electronic check,39.7,710.05,0,19,59,0.0,4034,0,Mount Shasta,0,0,Fiber Optic,41.33832,-122.290756,0,39.7,0,0,None,7309,0,0,0,1,19,0,0.0,0.0,0.0,710.05,1,1,96067
3244,1,0,0,0,10,1,1,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),54.5,568.2,0,29,59,33.98,4163,0,Nubieber,0,1,Fiber Optic,41.082471999999996,-121.19521499999999,0,54.5,0,0,None,240,0,0,0,0,10,0,0.0,339.7999999999999,0.0,568.2,1,1,96068
3245,0,0,1,1,23,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,83.8,1900.25,1,45,31,38.81,5737,1,Oak Run,1,0,DSL,40.689243,-122.037023,1,87.152,0,0,None,829,1,0,0,0,23,2,0.0,892.6300000000001,0.0,1900.25,0,1,96069
3246,1,0,0,0,3,1,0,DSL,0,0,1,0,Month-to-month,0,Mailed check,55.15,159.15,1,25,56,22.77,5698,1,Old Station,0,1,DSL,40.656287,-121.42896499999999,0,57.356,0,0,Offer E,182,0,2,0,1,3,2,0.0,68.31,0.0,159.15,1,1,96071
3247,0,0,0,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),111.6,8012.75,0,42,13,24.19,5425,0,Palo Cedro,1,0,DSL,40.582399,-122.19551200000001,0,111.6,0,0,None,4931,1,1,0,1,72,1,104.17,1741.68,0.0,8012.75,0,1,96073
3248,1,1,1,0,10,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.65,856.65,1,74,4,46.5,4990,1,Paskenta,0,1,Fiber Optic,39.884395,-122.58751299999999,1,90.116,0,2,None,263,0,2,1,0,10,3,0.0,465.0,0.0,856.65,0,1,96074
3249,0,0,1,1,10,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,55.55,551.3,0,30,59,5.74,2530,0,Paynes Creek,1,0,Cable,40.343213,-121.81541200000001,1,55.55,2,6,None,433,0,0,1,0,10,2,32.53,57.40000000000001,0.0,551.3,0,1,96075
3250,1,0,1,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.55,184.95,0,34,0,26.11,3971,0,Platina,0,1,NA,40.367964,-122.937379,1,20.55,0,6,None,215,0,2,1,0,11,2,0.0,287.21,0.0,184.95,0,0,96076
3251,0,1,0,0,37,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),106.75,4056.75,1,77,2,41.85,5849,1,Red Bluff,0,0,Fiber Optic,40.186772,-122.388361,0,111.02,0,0,Offer C,26438,0,0,0,0,37,5,81.0,1548.45,0.0,4056.75,0,0,96080
3252,1,0,1,1,17,1,1,DSL,1,0,0,0,One year,1,Mailed check,62.1,1096.65,0,58,28,32.27,3937,0,Round Mountain,0,1,Fiber Optic,40.923558,-122.059933,1,62.1,3,10,None,459,1,0,1,0,17,1,307.0,548.59,0.0,1096.65,0,0,96084
3253,0,0,1,1,36,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Credit card (automatic),104.5,3684.95,0,39,26,43.7,4102,0,Scott Bar,1,0,Fiber Optic,41.737961999999996,-123.07557,1,104.5,1,4,None,88,0,2,1,1,36,1,958.0,1573.2,0.0,3684.95,0,0,96085
3254,1,1,0,0,17,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.8,1752.45,0,77,25,17.26,3296,0,Seiad Valley,1,1,Fiber Optic,41.924174,-123.26078799999999,0,101.8,0,0,None,332,0,0,0,0,17,0,0.0,293.42,27.15,1752.45,0,1,96086
3255,0,1,1,1,66,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),110.6,7210.85,0,70,28,44.38,5418,0,Shasta,0,0,Cable,40.617614,-122.51286100000002,1,110.6,2,1,None,528,1,1,1,0,66,2,0.0,2929.080000000001,0.0,7210.85,0,1,96087
3256,1,0,1,1,61,1,0,DSL,1,1,1,1,One year,0,Bank transfer (automatic),84.9,5264.5,0,21,48,12.72,4413,0,Shingletown,1,1,DSL,40.497440999999995,-121.827524,1,84.9,2,3,Offer B,4231,1,0,1,1,61,0,2527.0,775.9200000000002,0.0,5264.5,1,0,96088
3257,1,0,0,0,22,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Mailed check,93.2,2157.3,0,50,17,46.5,4093,0,Tehama,0,1,DSL,40.021786999999996,-122.127576,0,93.2,0,0,None,405,0,0,0,1,22,0,0.0,1023.0,0.0,2157.3,0,1,96090
3258,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.4,24.4,0,40,6,0.0,3145,0,Trinity Center,0,1,Fiber Optic,41.081846999999996,-122.70054499999999,0,24.4,0,0,Offer E,734,0,0,0,0,1,0,0.0,0.0,0.0,24.4,0,0,96091
3259,0,0,0,0,6,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),70.55,433.95,0,52,27,30.54,4059,0,Vina,0,0,DSL,39.955164,-122.01856699999999,0,70.55,0,0,Offer E,439,0,0,0,0,6,1,0.0,183.24,0.0,433.95,0,1,96092
3260,1,0,0,0,31,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,78.45,2435.15,1,46,22,34.38,3091,1,Weaverville,0,1,Cable,40.759401000000004,-122.93933700000001,0,81.58800000000002,0,0,None,3749,1,1,0,0,31,3,536.0,1065.78,0.0,2435.15,0,0,96093
3261,0,0,1,1,68,1,0,DSL,1,1,1,1,Two year,1,Credit card (automatic),85.0,5607.75,0,61,16,6.28,6221,0,Weed,1,0,Cable,41.465121,-122.38094699999999,1,85.0,1,7,None,5896,1,0,1,1,68,2,0.0,427.04,0.0,5607.75,0,1,96094
3262,0,0,1,1,34,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,87.45,2874.15,1,39,4,40.78,3358,1,Whitmore,1,0,DSL,40.637105,-121.906949,1,90.948,0,1,None,843,0,0,1,0,34,1,115.0,1386.52,0.0,2874.15,0,0,96096
3263,0,0,1,1,52,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),85.8,4433.3,0,61,24,16.87,5494,0,Yreka,1,0,Fiber Optic,41.764869,-122.67131599999999,1,85.8,1,3,Offer B,9538,1,0,1,0,52,1,0.0,877.24,0.0,4433.3,0,1,96097
3264,0,0,0,1,10,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,91.1,964.35,0,43,52,42.93,3857,0,Alturas,1,0,Fiber Optic,41.468877,-120.54229,0,91.1,3,0,None,5096,1,0,0,0,10,2,501.0,429.3,0.0,964.35,0,0,96101
3265,1,0,1,1,29,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.75,1974.8,1,36,18,11.24,2663,1,Blairsden Graeagle,0,1,Cable,39.783747,-120.661032,1,73.58,0,1,None,1839,0,0,1,0,29,5,0.0,325.96,0.0,1974.8,0,1,96103
3266,0,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.1,1460.85,0,39,0,14.17,4598,0,Cedarville,0,0,NA,41.505916,-120.152505,1,20.1,2,10,None,857,0,0,1,0,72,1,0.0,1020.24,0.0,1460.85,0,0,96104
3267,1,0,1,1,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.05,951.55,0,28,0,6.51,5183,0,Chilcoot,0,1,NA,39.872961,-120.198876,1,20.05,1,9,Offer B,650,0,0,1,0,47,0,0.0,305.97,0.0,951.55,1,0,96105
3268,1,0,1,1,24,1,1,DSL,1,0,1,1,One year,0,Mailed check,74.8,1821.2,0,57,10,8.67,5535,0,Clio,0,1,Fiber Optic,39.745805,-120.580882,1,74.8,1,9,None,88,0,0,1,1,24,1,182.0,208.08,0.0,1821.2,0,0,96106
3269,1,0,0,0,65,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),24.8,1600.95,0,50,0,45.87,5826,0,Coleville,0,1,NA,38.42528,-119.47574099999999,0,24.8,0,0,Offer B,1332,0,1,0,0,65,1,0.0,2981.55,0.0,1600.95,0,0,96107
3270,0,0,0,0,4,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,100.85,399.25,0,31,3,7.94,5354,0,Davis Creek,0,0,DSL,41.750353999999994,-120.403885,0,100.85,0,0,Offer E,104,1,0,0,1,4,1,12.0,31.76,0.0,399.25,0,0,96108
3271,1,1,1,0,12,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.35,1218.55,1,66,4,48.5,3967,1,Doyle,0,1,Fiber Optic,40.012675,-120.10185700000001,1,105.404,0,1,None,1177,0,2,1,0,12,1,49.0,582.0,0.0,1218.55,0,0,96109
3272,1,0,0,0,1,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,81.7,81.7,1,31,31,9.81,5574,1,Eagleville,0,1,DSL,41.280341,-120.15038100000001,0,84.96799999999999,0,0,Offer E,132,0,2,0,0,1,5,0.0,9.81,0.0,81.7,0,0,96110
3273,1,0,0,0,33,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,68.25,2171.15,1,37,25,28.84,5647,1,Fort Bidwell,0,1,DSL,41.932207,-120.13594099999999,0,70.98,0,0,None,231,0,2,0,0,33,6,0.0,951.72,0.0,2171.15,0,1,96112
3274,0,0,0,0,34,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.1,3634.8,0,38,2,2.82,3941,0,Herlong,1,0,DSL,40.198234,-120.18088999999999,0,105.1,0,0,None,946,1,0,0,1,34,1,0.0,95.88,0.0,3634.8,0,1,96113
3275,0,0,1,0,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.4,292.4,0,46,0,14.61,4556,0,Janesville,0,0,NA,40.294034,-120.512622,1,20.4,0,0,None,3093,0,0,0,0,14,0,0.0,204.54,0.0,292.4,0,0,96114
3276,0,0,0,0,4,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.15,317.25,1,41,25,36.91,5762,1,Fallbrook,0,0,Cable,33.362575,-117.299644,0,82.316,0,0,Offer E,42239,0,0,0,1,4,1,0.0,147.64,0.0,317.25,0,1,92028
3277,1,0,1,1,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.0,218.55,0,54,0,4.26,5651,0,Likely,0,1,NA,41.266008,-120.49073100000001,1,20.0,2,7,None,277,0,0,1,0,13,0,0.0,55.38,0.0,218.55,0,0,96116
3278,0,0,1,1,65,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),79.4,5071.9,0,42,13,1.83,4023,0,Litchfield,0,0,Cable,40.507272,-120.338228,1,79.4,1,10,Offer B,385,1,0,1,1,65,1,0.0,118.95,0.0,5071.9,0,1,96117
3279,1,0,1,1,23,1,0,DSL,1,0,0,0,One year,0,Credit card (automatic),57.2,1423.35,0,59,30,37.86,4021,0,Loyalton,0,1,Fiber Optic,39.637471000000005,-120.22633799999998,1,57.2,2,4,None,1822,1,0,1,0,23,0,427.0,870.78,0.0,1423.35,0,0,96118
3280,1,0,1,0,55,1,0,DSL,1,1,0,0,Two year,0,Electronic check,58.6,3068.6,0,38,23,6.63,6231,0,Madeline,1,1,Cable,41.042003,-120.50608600000001,1,58.6,0,9,Offer B,85,0,0,1,0,55,0,0.0,364.65,0.0,3068.6,0,1,96119
3281,1,0,1,0,49,1,0,Fiber optic,0,1,1,1,Two year,1,Electronic check,94.8,4690.65,0,58,9,36.3,4252,0,Markleeville,0,1,DSL,38.735789000000004,-119.85798,1,94.8,0,8,Offer B,957,0,0,1,1,49,1,0.0,1778.6999999999996,0.0,4690.65,0,1,96120
3282,1,0,1,0,60,1,1,Fiber optic,0,1,1,1,One year,0,Bank transfer (automatic),102.5,6157.6,0,48,4,19.22,4968,0,Milford,1,1,DSL,40.181278999999996,-120.392967,1,102.5,0,8,Offer B,481,0,0,1,1,60,1,246.0,1153.1999999999996,0.0,6157.6,0,0,96121
3283,0,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.35,1442.65,0,24,0,23.47,5188,0,Portola,0,0,NA,39.786755,-120.445626,1,20.35,2,5,None,4236,0,0,1,0,69,0,0.0,1619.4299999999996,0.0,1442.65,1,0,96122
3284,1,0,0,0,40,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.9,3369.05,0,59,27,17.83,2904,0,Ravendale,0,1,Cable,40.845738,-120.32221899999999,0,84.9,0,0,None,61,0,0,0,0,40,0,910.0,713.1999999999998,0.0,3369.05,0,0,96123
3285,1,0,1,0,67,1,0,DSL,1,1,0,1,Two year,1,Credit card (automatic),69.2,4671.65,0,59,20,47.46,4323,0,Calpine,0,1,Fiber Optic,39.672813,-120.456699,1,69.2,0,0,None,322,1,0,0,1,67,2,0.0,3179.82,0.0,4671.65,0,1,96124
3286,1,1,0,0,35,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.45,3474.05,1,70,32,35.1,2080,1,Sierra City,0,1,DSL,39.600599,-120.636358,0,99.26799999999999,0,0,Offer C,348,0,0,0,0,35,0,1112.0,1228.5,0.0,3474.05,0,0,96125
3287,1,0,1,1,19,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,100.95,1875.55,1,29,56,5.93,4072,1,Sierraville,0,1,DSL,39.559709000000005,-120.34563899999999,1,104.988,0,1,None,227,1,0,1,1,19,2,1050.0,112.67,0.0,1875.55,1,0,96126
3288,0,0,1,1,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.85,272.35,0,56,0,27.62,3163,0,Standish,0,0,NA,40.346634,-120.386422,1,20.85,3,6,None,408,0,1,1,0,13,1,0.0,359.06,0.0,272.35,0,0,96128
3289,0,0,0,1,41,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),88.5,3645.05,0,33,10,18.72,5984,0,Susanville,0,0,Fiber Optic,40.559177000000005,-120.612113,0,88.5,2,0,None,19440,0,0,0,0,41,0,365.0,767.52,0.0,3645.05,0,0,96130
3290,0,0,0,0,4,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,35.0,135.75,0,46,26,0.0,3523,0,Termo,1,0,Fiber Optic,41.027281,-120.669427,0,35.0,0,0,None,72,0,0,0,0,4,1,3.53,0.0,0.0,135.75,0,1,96132
3291,0,0,1,1,24,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,55.15,1319.85,0,29,85,27.37,2200,0,Topaz,0,0,Cable,38.636052,-119.48916200000001,1,55.15,3,7,None,116,1,0,1,0,24,3,1122.0,656.88,0.0,1319.85,1,0,96133
3292,0,0,0,0,5,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Credit card (automatic),50.95,229.4,0,46,26,0.0,3573,0,Tulelake,0,0,Fiber Optic,41.813521,-121.49266599999999,0,50.95,0,0,Offer E,2595,0,0,0,1,5,1,0.0,0.0,0.0,229.4,0,1,96134
3293,0,0,0,0,5,1,1,DSL,0,1,0,1,Month-to-month,1,Electronic check,64.0,370.25,0,37,29,44.78,4421,0,Wendel,0,0,DSL,40.345949,-120.08118700000001,0,64.0,0,0,None,162,0,0,0,1,5,1,0.0,223.9,0.0,370.25,0,1,96136
3294,0,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.1,69.1,1,46,21,16.55,4779,1,Westwood,0,0,Cable,40.271535,-121.01808700000001,1,71.86399999999998,0,1,Offer E,4158,0,0,1,0,1,0,0.0,16.55,0.0,69.1,0,0,96137
3295,0,0,1,1,72,1,1,DSL,1,1,1,0,Two year,0,Bank transfer (automatic),80.2,5714.2,0,39,23,49.12,6087,0,Carnelian Bay,1,0,Cable,39.227434,-120.091806,1,80.2,3,7,None,1943,1,0,1,0,72,0,1314.0,3536.64,0.0,5714.2,0,0,96140
3296,0,0,0,0,24,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),49.3,1233.25,0,34,16,4.82,5394,0,Homewood,1,0,DSL,39.117018,-120.212535,0,49.3,0,0,None,858,0,0,0,0,24,1,197.0,115.68,0.0,1233.25,0,0,96141
3297,0,0,1,0,42,1,1,DSL,1,0,1,1,Two year,0,Credit card (automatic),84.35,3571.6,0,25,52,9.84,3363,0,Tahoma,1,0,DSL,39.061227,-120.179546,1,84.35,0,4,None,1291,1,2,1,1,42,2,1857.0,413.28,0.0,3571.6,1,0,96142
3298,0,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,83.3,0,33,0,25.8,4596,0,Kings Beach,0,0,NA,39.246654,-120.029273,0,20.05,0,0,None,4806,0,0,0,0,4,0,0.0,103.2,0.0,83.3,0,0,96143
3299,1,0,0,0,68,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),117.2,8035.95,0,39,3,32.67,4629,0,Tahoe City,1,1,DSL,39.178337,-120.162806,0,117.2,0,0,None,4002,1,0,0,1,68,0,0.0,2221.56,0.0,8035.95,0,1,96145
3300,0,0,1,1,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,579.4,0,23,0,28.4,3342,0,Olympic Valley,0,0,NA,39.191796999999994,-120.212401,1,20.1,3,3,None,942,0,0,1,0,33,0,0.0,937.2,0.0,579.4,1,0,96146
3301,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.6,69.6,1,68,11,45.8,2151,1,Tahoe Vista,0,0,DSL,39.241240000000005,-120.05476499999999,0,72.384,0,0,Offer E,678,0,0,0,0,1,4,0.0,45.8,0.0,69.6,0,0,96148
3302,1,0,0,0,31,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,103.45,3066.45,1,53,33,9.27,5387,1,South Lake Tahoe,1,1,Fiber Optic,38.911577,-120.106169,0,107.588,0,0,None,33038,0,0,0,1,31,2,0.0,287.37,0.0,3066.45,0,1,96150
3303,0,0,0,0,4,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),77.95,305.55,1,31,29,30.95,5365,1,San Diego,0,0,DSL,32.957195,-117.202542,0,81.06800000000001,0,0,None,28201,0,1,0,0,4,2,89.0,123.8,0.0,305.55,0,0,92130
3304,1,1,1,0,69,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,109.95,7634.25,0,71,17,18.41,4297,0,Los Angeles,1,1,Cable,33.973616,-118.24902,1,109.95,0,1,None,54492,1,0,1,0,69,0,0.0,1270.29,0.0,7634.25,0,1,90001
3305,1,1,0,0,38,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,94.75,3653,0,68,13,46.96,3654,0,Los Angeles,0,1,Fiber Optic,33.949255,-118.246978,0,94.75,0,0,None,44586,0,0,0,0,38,0,0.0,1784.48,45.82,3653.0,0,1,90002
3306,0,0,1,1,3,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.0,241.3,0,49,22,19.18,4264,0,Los Angeles,0,0,Cable,33.964131,-118.272783,1,80.0,3,2,None,58198,1,0,1,0,3,0,53.0,57.54,0.0,241.3,0,0,90003
3307,0,0,1,1,48,1,1,DSL,0,1,1,1,Two year,0,Electronic check,79.65,3870.3,0,44,27,8.94,3246,0,Los Angeles,0,0,DSL,34.076259,-118.31071499999999,1,79.65,1,5,None,67852,1,0,1,1,48,0,0.0,429.12,0.0,3870.3,0,1,90004
3308,0,0,1,0,15,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.2,387.9,0,35,0,46.68,4411,0,Los Angeles,0,0,NA,34.059281,-118.30742,1,25.2,0,9,None,43019,0,0,1,0,15,0,0.0,700.2,0.0,387.9,0,0,90005
3309,0,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.9,527.5,0,50,0,1.36,3048,0,Los Angeles,0,0,NA,34.048013,-118.293953,0,19.9,0,0,None,62784,0,0,0,0,25,1,0.0,34.0,0.0,527.5,0,0,90006
3310,0,1,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,78.45,78.45,1,65,14,18.37,2139,1,Los Angeles,0,0,Cable,34.027337,-118.28515,0,81.58800000000002,0,0,Offer E,45025,0,2,0,0,1,1,0.0,18.37,0.0,78.45,0,0,90007
3311,0,0,0,0,48,0,No phone service,DSL,1,1,1,0,Month-to-month,1,Electronic check,44.8,2104.55,0,62,23,0.0,2469,0,Los Angeles,0,0,DSL,34.008293,-118.34676599999999,0,44.8,0,0,None,30852,0,0,0,0,48,0,0.0,0.0,0.0,2104.55,0,1,90008
3312,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.3,20.3,0,29,0,10.84,4270,0,Los Angeles,0,1,NA,34.062125,-118.31570900000001,0,20.3,0,0,None,1957,0,1,0,0,1,2,0.0,10.84,0.0,20.3,1,0,90010
3313,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.2,19.2,0,22,0,26.37,2716,0,Los Angeles,0,1,NA,34.007090000000005,-118.25868100000001,0,19.2,0,0,None,101215,0,0,0,0,1,0,0.0,26.37,0.0,19.2,1,0,90011
3314,0,0,0,0,37,1,0,Fiber optic,0,1,0,0,One year,0,Electronic check,80.05,3019.1,0,48,11,9.61,3364,0,Los Angeles,1,0,Cable,34.065875,-118.23872800000001,0,80.05,0,0,None,30596,0,0,0,0,37,0,332.0,355.57,0.0,3019.1,0,0,90012
3315,1,1,1,0,66,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),107.35,7051.95,0,71,26,7.86,4138,0,Los Angeles,1,1,Fiber Optic,34.044639000000004,-118.24041299999999,1,107.35,0,7,None,9732,1,0,1,0,66,1,0.0,518.76,39.18,7051.95,0,1,90013
3316,0,0,1,0,26,0,No phone service,DSL,1,1,1,0,One year,0,Bank transfer (automatic),47.85,1190.5,0,34,28,0.0,4362,0,Los Angeles,1,0,Fiber Optic,34.043144,-118.251977,1,47.85,0,10,None,3524,0,0,1,0,26,2,0.0,0.0,0.0,1190.5,0,1,90014
3317,1,0,1,0,63,1,0,DSL,1,1,1,0,One year,0,Credit card (automatic),70.8,4448.8,0,59,13,46.99,5114,0,Los Angeles,0,1,DSL,34.039224,-118.26629299999999,1,70.8,0,6,None,15140,1,0,1,0,63,0,0.0,2960.370000000001,0.0,4448.8,0,1,90015
3318,1,0,0,0,10,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,29.5,255.25,1,46,33,0.0,3797,1,Los Angeles,1,1,Fiber Optic,34.028331,-118.35433799999998,0,30.68,0,0,Offer D,46984,0,0,0,0,10,0,84.0,0.0,0.0,255.25,0,0,90016
3319,0,0,0,0,2,1,0,DSL,1,0,1,1,Month-to-month,1,Electronic check,70.75,146.9,1,64,11,26.93,3257,1,Los Angeles,0,0,DSL,34.052842,-118.264495,0,73.58,0,0,None,20692,0,1,0,1,2,4,16.0,53.86,0.0,146.9,0,0,90017
3320,1,1,1,0,18,1,0,DSL,1,0,0,1,Month-to-month,1,Credit card (automatic),59.1,1011.05,0,74,13,5.73,2422,0,Los Angeles,0,1,Fiber Optic,34.028735,-118.31723600000001,1,59.1,0,6,None,47143,0,0,1,0,18,1,131.0,103.14,31.05,1011.05,0,0,90018
3321,0,0,1,0,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.55,1714.95,0,40,0,49.39,4312,0,Los Angeles,0,0,NA,34.049841,-118.33846000000001,1,25.55,0,9,None,67520,0,0,1,0,64,1,0.0,3160.96,0.0,1714.95,0,0,90019
3322,0,1,0,0,9,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.45,762.5,1,76,23,12.91,3543,1,San Diego,0,0,Fiber Optic,32.898613,-117.202937,0,87.82799999999999,0,0,Offer E,4258,0,0,0,0,9,3,175.0,116.19,0.0,762.5,0,0,92121
3323,0,0,0,1,28,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,535.35,0,27,0,26.09,4476,0,Los Angeles,0,0,NA,34.029043,-118.23950400000001,0,20.25,3,0,None,3012,0,0,0,0,28,0,0.0,730.52,0.0,535.35,1,0,90021
3324,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.55,75.55,0,32,26,7.11,3503,0,Los Angeles,1,0,Fiber Optic,34.02381,-118.156582,0,75.55,0,0,None,68701,0,0,0,0,1,1,0.0,7.11,0.0,75.55,0,0,90022
3325,1,0,0,0,4,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.65,338.9,1,19,58,6.91,2330,1,Los Angeles,0,1,Cable,34.017697,-118.200577,0,89.07600000000002,0,0,None,47487,0,3,0,1,4,2,0.0,27.64,0.0,338.9,1,1,90023
3326,1,1,0,0,38,1,0,DSL,0,1,1,0,One year,1,Credit card (automatic),70.15,2497.35,1,73,33,5.75,2645,1,Los Angeles,1,1,DSL,34.066303000000005,-118.435479,0,72.956,0,0,Offer C,44150,1,2,0,0,38,2,824.0,218.5,0.0,2497.35,0,0,90024
3327,1,0,1,0,66,1,1,Fiber optic,0,1,0,1,One year,0,Electronic check,95.3,6273.4,0,36,24,25.83,5706,0,Los Angeles,1,1,Fiber Optic,34.046174,-118.44633300000001,1,95.3,0,1,None,41175,0,0,1,1,66,0,150.56,1704.78,0.0,6273.4,0,1,90025
3328,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.25,70.25,0,20,51,10.05,4063,0,Los Angeles,0,0,Fiber Optic,34.078990999999995,-118.26380400000001,0,70.25,0,0,None,73686,0,1,0,0,1,1,0.0,10.05,0.0,70.25,1,1,90026
3329,0,0,1,0,18,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.3,908.75,0,42,17,35.96,3740,0,Los Angeles,0,0,Fiber Optic,34.127194,-118.295647,1,50.3,0,4,Offer D,48727,1,0,1,0,18,1,0.0,647.28,0.0,908.75,0,1,90027
3330,1,1,0,0,51,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,97.8,4913.3,1,70,12,19.49,6204,1,Los Angeles,1,1,Fiber Optic,34.099869,-118.326843,0,101.712,0,0,Offer B,30568,0,0,0,0,51,1,0.0,993.99,0.0,4913.3,0,1,90028
3331,1,0,1,1,0,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.85, ,0,56,0,15.51,2019,0,Los Angeles,0,1,NA,34.089953,-118.294824,1,19.85,1,5,None,41713,0,0,1,0,10,2,0.0,155.1,0.0,198.5,0,0,90029
3332,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,46.3,46.3,1,39,23,48.22,3017,1,Los Angeles,0,1,Cable,34.085807,-118.206617,0,48.152,0,0,None,38415,0,1,0,0,1,3,0.0,48.22,0.0,46.3,0,0,90031
3333,1,0,0,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.35,212.3,0,44,0,17.23,2558,0,Los Angeles,0,1,NA,34.078821000000005,-118.177576,0,19.35,3,0,Offer D,46960,0,0,0,0,12,1,0.0,206.76,0.0,212.3,0,0,90032
3334,0,0,0,0,41,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.3,4443.45,1,63,24,10.43,5383,1,Los Angeles,1,0,Fiber Optic,34.050197999999995,-118.21094599999999,0,110.552,0,0,None,49431,0,0,0,1,41,0,1066.0,427.63,0.0,4443.45,0,0,90033
3335,1,0,0,0,12,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,25.0,316.2,0,37,0,2.29,4408,0,Los Angeles,0,1,NA,34.030578000000006,-118.39961299999999,0,25.0,0,0,Offer D,58218,0,0,0,0,12,0,0.0,27.48,0.0,316.2,0,0,90034
3336,0,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.3,1079.05,0,62,0,3.18,5153,0,Los Angeles,0,0,NA,34.051809000000006,-118.383843,1,20.3,1,3,None,27799,0,0,1,0,55,0,0.0,174.9,0.0,1079.05,0,0,90035
3337,0,0,0,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.35,564.65,0,63,17,25.17,4989,0,Los Angeles,0,0,DSL,34.070291,-118.34919099999999,0,75.35,0,0,None,32901,0,0,0,0,7,2,96.0,176.19,0.0,564.65,0,0,90036
3338,0,0,0,0,12,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.4,1095.65,1,36,10,17.46,5047,1,Los Angeles,1,0,Cable,34.002642,-118.287596,0,92.976,0,0,Offer D,56709,1,2,0,1,12,3,0.0,209.52,0.0,1095.65,0,1,90037
3339,0,0,1,1,68,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),88.0,6161.9,0,49,22,43.51,5436,0,Los Angeles,1,0,DSL,34.088017,-118.327168,1,88.0,1,10,None,32562,1,0,1,1,68,0,1356.0,2958.68,0.0,6161.9,0,0,90038
3340,0,1,0,0,5,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),83.15,446.05,1,68,28,41.83,2516,1,Los Angeles,0,0,DSL,34.110845,-118.25959499999999,0,86.47600000000001,0,0,None,29310,0,1,0,0,5,2,125.0,209.15,0.0,446.05,0,0,90039
3341,0,1,0,0,49,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,43.8,2106.05,0,78,3,35.65,5651,0,Los Angeles,0,0,DSL,33.994524,-118.149953,0,43.8,0,0,None,9805,0,0,0,0,49,2,0.0,1746.85,20.45,2106.05,0,1,90040
3342,1,0,0,0,40,0,No phone service,DSL,1,1,1,1,One year,0,Credit card (automatic),62.05,2511.55,0,38,19,0.0,2290,0,Los Angeles,1,1,Cable,34.137412,-118.20760700000001,0,62.05,0,0,None,27866,0,0,0,1,40,0,0.0,0.0,0.0,2511.55,0,1,90041
3343,0,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.1,318.6,0,23,0,47.25,4545,0,Los Angeles,0,0,NA,34.11572,-118.19275400000001,0,20.1,0,0,Offer D,64672,0,0,0,0,16,0,0.0,756.0,0.0,318.6,1,0,90042
3344,1,0,0,0,10,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.15,811.8,1,28,94,29.24,4231,1,Los Angeles,0,1,DSL,33.988543,-118.33408100000001,0,77.11600000000001,0,0,Offer D,44764,0,0,0,1,10,7,763.0,292.4,0.0,811.8,1,0,90043
3345,0,0,1,0,72,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,101.35,7323.15,0,49,23,46.1,4497,0,Los Angeles,1,0,Fiber Optic,33.952714,-118.292061,1,101.35,0,6,Offer A,87383,0,0,1,1,72,0,168.43,3319.2000000000007,0.0,7323.15,0,1,90044
3346,0,1,0,0,2,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.05,186.05,0,70,22,21.9,5039,0,Los Angeles,0,0,Fiber Optic,33.954017,-118.402447,0,84.05,0,0,Offer E,39334,0,0,0,0,2,0,41.0,43.8,0.0,186.05,0,0,90045
3347,1,0,1,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.9,454,0,32,0,18.91,4076,0,Los Angeles,0,1,NA,34.108455,-118.362081,1,20.9,1,1,Offer D,49839,0,1,1,0,23,1,0.0,434.93,0.0,454.0,0,0,90046
3348,0,1,0,0,71,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,105.9,7521.95,0,65,23,25.61,5479,0,Los Angeles,1,0,DSL,33.958149,-118.30844099999999,0,105.9,0,0,None,47107,0,0,0,1,71,2,0.0,1818.31,6.65,7521.95,0,1,90047
3349,0,0,1,0,11,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.5,1056.95,1,43,29,31.08,5286,1,Los Angeles,1,0,Cable,34.072945000000004,-118.37267,1,103.48,0,1,Offer D,21739,0,1,1,1,11,2,0.0,341.88,0.0,1056.95,0,1,90048
3350,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.15,44.15,1,44,11,8.77,4773,1,Los Angeles,0,1,Cable,34.091829,-118.491244,0,45.916000000000004,0,0,None,33523,0,0,0,0,1,1,0.0,8.77,0.0,44.15,0,0,90049
3351,0,0,0,0,16,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,53.9,834.15,1,36,9,6.86,5091,1,Los Angeles,0,0,Fiber Optic,33.987945,-118.370442,0,56.056000000000004,0,0,Offer D,8115,1,0,0,0,16,6,75.0,109.76,0.0,834.15,0,0,90056
3352,0,0,0,0,1,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Mailed check,85.45,85.45,1,22,30,31.03,2318,1,Los Angeles,0,0,Fiber Optic,34.061918,-118.27793899999999,0,88.86800000000002,0,0,None,44004,0,0,0,1,1,4,0.0,31.03,0.0,85.45,1,1,90057
3353,1,0,1,0,12,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),85.05,999.8,0,44,20,44.6,2540,0,Los Angeles,0,1,Fiber Optic,34.001616999999996,-118.222274,1,85.05,0,1,Offer D,3642,0,0,1,1,12,3,0.0,535.2,0.0,999.8,0,1,90058
3354,0,0,0,0,54,0,No phone service,DSL,1,0,0,1,One year,0,Bank transfer (automatic),44.1,2369.7,0,52,21,0.0,6205,0,Los Angeles,0,0,Fiber Optic,33.927254,-118.249826,0,44.1,0,0,None,38128,1,0,0,1,54,1,0.0,0.0,0.0,2369.7,0,1,90059
3355,0,0,1,0,68,1,1,Fiber optic,0,1,0,0,Two year,0,Credit card (automatic),90.2,6297.65,0,27,26,3.41,4095,0,Los Angeles,1,0,Cable,33.921279999999996,-118.27418600000001,1,90.2,0,3,Offer A,24511,1,0,1,0,68,0,0.0,231.88,0.0,6297.65,1,1,90061
3356,0,0,1,1,4,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.85,239.55,1,36,24,12.88,5386,1,Los Angeles,0,0,Cable,34.003553000000004,-118.30893300000001,1,52.88399999999999,1,1,None,29299,0,1,1,0,4,2,57.0,51.52,0.0,239.55,0,0,90062
3357,0,0,0,1,1,1,0,DSL,0,0,0,1,Month-to-month,0,Electronic check,59.2,59.2,1,40,26,13.58,5020,1,Los Angeles,1,0,Cable,34.044271,-118.18523700000001,0,61.56800000000001,3,0,None,55668,0,1,0,1,1,7,0.0,13.58,0.0,59.2,0,0,90063
3358,1,0,0,0,27,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,53.45,1461.45,0,53,28,15.09,2191,0,Los Angeles,0,1,DSL,34.037251,-118.423573,0,53.45,0,0,None,24505,1,1,0,0,27,1,409.0,407.43,0.0,1461.45,0,0,90064
3359,1,0,0,0,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.95,416.4,0,34,0,44.01,3632,0,Los Angeles,0,1,NA,34.108833000000004,-118.22971499999998,0,19.95,0,0,Offer D,47534,0,0,0,0,21,0,0.0,924.21,0.0,416.4,0,0,90065
3360,1,0,0,0,13,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,83.2,1060.6,1,42,20,35.4,4028,1,Los Angeles,1,1,Fiber Optic,34.002028,-118.430656,0,86.52799999999999,0,0,Offer D,55204,0,0,0,0,13,3,0.0,460.2,0.0,1060.6,0,1,90066
3361,0,1,0,0,64,1,1,DSL,0,1,0,1,Month-to-month,0,Credit card (automatic),74.65,4869.35,0,68,21,27.7,5113,0,Los Angeles,1,0,Fiber Optic,34.057496,-118.413959,0,74.65,0,0,None,2527,1,0,0,0,64,1,0.0,1772.8,47.04,4869.35,0,1,90067
3362,0,0,0,0,1,1,0,DSL,1,1,0,0,Month-to-month,1,Electronic check,54.9,54.9,1,19,64,44.36,2833,1,Los Angeles,0,0,DSL,34.137411,-118.328915,0,57.096,0,0,None,21728,0,3,0,1,1,2,0.0,44.36,0.0,54.9,1,0,90068
3363,1,0,1,0,57,0,No phone service,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),57.5,3265.95,0,27,69,0.0,4133,0,West Hollywood,1,1,DSL,34.093781,-118.38106100000002,1,57.5,0,2,None,20408,1,0,1,1,57,2,0.0,0.0,0.0,3265.95,1,1,90069
3364,0,0,1,0,21,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,103.9,2254.2,1,57,18,1.21,3769,1,Los Angeles,1,0,Cable,34.052917,-118.255178,1,108.056,0,1,Offer D,21,0,0,1,1,21,1,0.0,25.41,0.0,2254.2,0,1,90071
3365,1,0,0,0,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.65,358.15,0,25,0,34.68,5596,0,Los Angeles,0,1,NA,34.102084000000005,-118.451629,0,19.65,0,0,Offer D,10470,0,0,0,0,19,0,0.0,658.92,0.0,358.15,1,0,90077
3366,1,0,1,0,31,1,0,Fiber optic,0,0,1,1,One year,1,Electronic check,93.8,2939.8,0,27,52,36.69,2510,0,Bell,1,1,DSL,33.970343,-118.17136799999999,1,93.8,0,2,None,105285,0,0,1,1,31,0,0.0,1137.39,0.0,2939.8,1,1,90201
3367,1,0,0,0,52,1,1,DSL,1,1,1,1,Two year,1,Mailed check,89.25,4652.4,0,34,30,6.8,4624,0,Beverly Hills,1,1,DSL,34.099891,-118.41433799999999,0,89.25,0,0,None,21397,1,0,0,1,52,1,1396.0,353.6,0.0,4652.4,0,0,90210
3368,0,0,0,0,46,1,1,Fiber optic,0,1,0,1,One year,1,Electronic check,94.15,4408.45,0,55,3,33.18,3924,0,Beverly Hills,1,0,DSL,34.063947,-118.38300100000001,0,94.15,0,0,None,8321,0,0,0,1,46,0,13.23,1526.28,0.0,4408.45,0,1,90211
3369,0,1,0,0,11,1,1,DSL,1,0,0,0,Month-to-month,1,Electronic check,55.6,580.8,0,73,3,2.81,5014,0,Beverly Hills,0,0,Cable,34.062095,-118.401508,0,55.6,0,0,None,11355,0,0,0,0,11,0,17.0,30.91,15.2,580.8,0,0,90212
3370,0,0,1,1,53,0,No phone service,DSL,1,1,0,1,Month-to-month,1,Bank transfer (automatic),48.7,2495.2,0,40,25,0.0,4116,0,Compton,1,0,DSL,33.88151,-118.234451,1,48.7,3,5,None,47305,0,0,1,1,53,1,0.0,0.0,0.0,2495.2,0,1,90220
3371,0,0,1,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.25,180.3,1,35,0,29.01,5638,1,Compton,0,0,NA,33.885811,-118.20645900000001,1,19.25,3,1,Offer D,51387,0,0,1,0,11,2,0.0,319.11,0.0,180.3,0,0,90221
3372,1,1,0,0,57,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),104.9,5913.95,0,68,15,32.12,5838,0,Compton,0,1,Fiber Optic,33.912246,-118.236773,0,104.9,0,0,None,29825,1,0,0,0,57,1,0.0,1830.84,1.69,5913.95,0,1,90222
3373,0,1,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,75.45,158.4,1,77,28,23.46,3350,1,Culver City,0,0,DSL,33.993990999999994,-118.39703999999999,0,78.468,0,0,None,31963,0,0,0,0,2,2,44.0,46.92,0.0,158.4,0,0,90230
3374,0,1,0,0,2,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,54.85,104.2,1,73,7,25.74,3016,1,Culver City,0,0,Cable,34.019323,-118.391902,0,57.044,0,0,None,15195,0,0,0,0,2,0,0.0,51.48,0.0,104.2,0,1,90232
3375,0,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.9,1389.35,0,34,0,12.22,5789,0,Downey,0,0,NA,33.956228,-118.120993,1,19.9,1,4,Offer A,24908,0,0,1,0,71,0,0.0,867.62,0.0,1389.35,0,0,90240
3376,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.4,19.4,0,58,0,48.79,3160,0,Downey,0,0,NA,33.940884000000004,-118.128628,1,19.4,2,6,None,40152,0,0,1,0,1,0,0.0,48.79,0.0,19.4,0,0,90241
3377,1,0,1,0,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.05,1629.2,0,19,0,25.19,4187,0,Downey,0,1,NA,33.921793,-118.140588,1,25.05,0,4,Offer A,42459,0,0,1,0,68,1,0.0,1712.92,0.0,1629.2,1,0,90242
3378,1,0,1,0,72,1,0,DSL,1,1,1,1,Two year,0,Mailed check,84.45,6033.1,0,35,26,35.06,6297,0,El Segundo,1,1,Cable,33.917145,-118.401554,1,84.45,0,8,Offer A,16041,1,0,1,1,72,1,0.0,2524.32,0.0,6033.1,0,1,90245
3379,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.3,44.4,0,34,0,49.91,3009,0,Gardena,0,0,NA,33.890853,-118.29796699999999,0,19.3,0,0,None,47758,0,1,0,0,2,1,0.0,99.82,0.0,44.4,0,0,90247
3380,1,1,1,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.1,95.1,1,71,12,4.89,5795,1,Gardena,0,1,Fiber Optic,33.876482,-118.284077,1,98.904,0,1,None,9960,0,0,1,0,1,6,0.0,4.89,0.0,95.1,0,1,90248
3381,0,0,0,0,41,1,0,DSL,1,0,1,1,One year,1,Bank transfer (automatic),79.85,3320.75,0,57,5,38.21,5556,0,Gardena,1,0,DSL,33.90139,-118.315697,0,79.85,0,0,None,26442,1,0,0,1,41,0,0.0,1566.61,0.0,3320.75,0,1,90249
3382,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.55,1867.7,0,53,0,36.82,6425,0,Hawthorne,0,1,NA,33.914775,-118.348083,1,25.55,3,4,Offer A,93315,0,0,1,0,72,2,0.0,2651.04,0.0,1867.7,0,0,90250
3383,1,0,1,0,6,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.5,438,1,33,14,21.23,5838,1,Hermosa Beach,0,1,Cable,33.865320000000004,-118.396336,1,78.52,0,4,None,18693,0,3,1,0,6,4,61.0,127.38,0.0,438.0,0,0,90254
3384,0,0,1,1,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.75,325.45,1,25,64,48.48,5026,1,Huntington Park,1,0,Cable,33.97803,-118.217141,1,76.7,0,5,None,78114,0,3,1,1,4,2,208.0,193.92,0.0,325.45,1,0,90255
3385,1,0,0,0,12,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.05,1148.1,1,39,28,44.71,2577,1,Lawndale,0,1,DSL,33.88856,-118.35181299999999,0,99.89200000000001,0,0,Offer D,33300,0,0,0,1,12,3,321.0,536.52,0.0,1148.1,0,0,90260
3386,0,0,1,0,58,1,1,DSL,1,0,0,1,One year,1,Electronic check,68.4,3972.25,0,24,53,26.99,5269,0,Lynwood,0,0,Fiber Optic,33.923573,-118.20066899999999,1,68.4,0,8,None,69850,1,0,1,1,58,1,0.0,1565.4199999999996,0.0,3972.25,1,1,90262
3387,0,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.65,155.9,0,55,0,15.54,2100,0,Malibu,0,0,NA,34.037037,-118.705803,0,20.65,0,0,None,11,0,0,0,0,7,1,0.0,108.78,0.0,155.9,0,0,90263
3388,0,0,1,0,65,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,55.15,3673.15,0,63,26,19.99,6205,0,Malibu,1,0,Fiber Optic,34.074571999999996,-118.831181,1,55.15,0,7,None,19630,0,1,1,0,65,3,95.5,1299.35,0.0,3673.15,0,1,90265
3389,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.6,70.6,0,31,14,36.12,3530,0,Manhattan Beach,0,1,Fiber Optic,33.889632,-118.39737,0,70.6,0,0,None,33758,0,0,0,0,1,0,0.0,36.12,0.0,70.6,0,0,90266
3390,1,0,1,0,56,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.95,1126.75,0,29,0,48.87,4838,0,Maywood,0,1,NA,33.988572,-118.18656499999999,1,19.95,0,0,None,28094,0,0,0,0,56,2,0.0,2736.72,0.0,1126.75,1,0,90270
3391,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.0,73.45,0,21,0,8.38,4345,0,Pacific Palisades,0,1,NA,34.079449,-118.54830600000001,0,19.0,0,0,None,22548,0,0,0,0,4,0,0.0,33.52,0.0,73.45,1,0,90272
3392,0,0,1,1,58,1,0,DSL,0,0,0,0,One year,1,Mailed check,44.1,2413.05,0,44,25,22.65,5040,0,Palos Verdes Peninsula,0,0,DSL,33.788208000000004,-118.404955,1,44.1,3,7,None,24979,0,0,1,0,58,0,603.0,1313.6999999999996,0.0,2413.05,0,0,90274
3393,1,0,1,0,62,1,1,Fiber optic,0,0,1,1,Two year,1,Bank transfer (automatic),107.6,6912.7,0,54,28,34.62,4697,0,Rancho Palos Verdes,1,1,Cable,33.753146,-118.36745900000001,1,107.6,0,8,None,41263,1,1,1,1,62,1,1936.0,2146.44,0.0,6912.7,0,0,90275
3394,1,0,0,0,26,1,1,DSL,1,1,0,0,One year,0,Electronic check,61.55,1581.95,0,23,73,38.04,5156,0,Redondo Beach,0,1,Fiber Optic,33.830453000000006,-118.384565,0,61.55,0,0,None,34191,0,0,0,0,26,0,1155.0,989.04,0.0,1581.95,1,0,90277
3395,1,0,0,0,62,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Bank transfer (automatic),90.7,5586.45,0,44,2,18.9,5496,0,Redondo Beach,1,1,Fiber Optic,33.873395,-118.37019,0,90.7,0,0,None,37322,0,0,0,0,62,2,0.0,1171.8,0.0,5586.45,0,1,90278
3396,0,0,1,1,58,1,0,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),99.25,5846.65,0,20,76,39.05,4098,0,South Gate,0,0,Fiber Optic,33.944624,-118.19261499999999,1,99.25,2,9,None,96267,0,0,1,1,58,1,0.0,2264.9,0.0,5846.65,1,1,90280
3397,0,0,1,0,68,1,1,DSL,1,1,1,1,Two year,1,Electronic check,91.7,6424.7,0,45,5,15.65,4113,0,Topanga,1,0,DSL,34.115192,-118.61017,1,91.7,0,10,Offer A,5451,1,0,1,1,68,1,32.12,1064.2,0.0,6424.7,0,1,90290
3398,0,0,1,1,61,1,1,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),100.7,6018.65,0,60,19,18.26,4804,0,Venice,1,0,Fiber Optic,33.991782,-118.479229,1,100.7,1,5,Offer B,31021,0,0,1,1,61,3,0.0,1113.86,0.0,6018.65,0,1,90291
3399,0,0,0,0,42,1,1,DSL,0,0,1,1,Two year,1,Credit card (automatic),78.45,3373.4,0,56,15,20.27,3192,0,Marina Del Rey,1,0,Fiber Optic,33.977468,-118.445475,0,78.45,0,0,Offer B,18058,1,0,0,1,42,1,506.0,851.34,0.0,3373.4,0,0,90292
3400,1,0,0,0,18,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Bank transfer (automatic),84.3,1537.9,0,19,73,2.26,4612,0,Playa Del Rey,0,1,DSL,33.947305,-118.43984099999999,0,84.3,0,0,Offer D,11264,0,0,0,0,18,0,1123.0,40.67999999999999,0.0,1537.9,1,0,90293
3401,0,0,0,0,56,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.55,1080.55,0,57,0,13.89,5764,0,Inglewood,0,0,NA,33.956445,-118.35863400000001,0,19.55,0,0,Offer B,37527,0,0,0,0,56,1,0.0,777.84,0.0,1080.55,0,0,90301
3402,0,0,0,0,4,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,88.95,355.2,1,30,56,48.32,5948,1,Inglewood,0,0,Cable,33.975332,-118.35525200000001,0,92.508,0,0,None,30779,0,4,0,1,4,2,0.0,193.28,0.0,355.2,0,1,90302
3403,0,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.45,82.85,0,31,0,3.05,4344,0,Inglewood,0,0,NA,33.936291,-118.33263899999999,0,20.45,0,0,None,27778,0,0,0,0,4,1,0.0,12.2,0.0,82.85,0,0,90303
3404,0,0,0,1,35,1,0,DSL,1,1,0,0,One year,0,Credit card (automatic),55.6,2016.45,0,46,56,12.56,5964,0,Inglewood,0,0,DSL,33.936827,-118.359824,0,55.6,3,0,None,28680,0,0,0,0,35,0,1129.0,439.6,0.0,2016.45,0,0,90304
3405,0,0,1,1,64,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),86.8,5327.25,0,31,12,27.74,4915,0,Inglewood,0,0,DSL,33.958134,-118.330905,1,86.8,2,0,Offer B,13779,1,0,0,0,64,0,639.0,1775.36,0.0,5327.25,0,0,90305
3406,0,0,0,0,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.95,683.25,0,23,0,31.79,5772,0,Santa Monica,0,0,NA,34.015481,-118.49323100000001,0,20.95,0,0,None,5221,0,0,0,0,31,1,0.0,985.49,0.0,683.25,1,0,90401
3407,0,1,1,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.05,1263.05,0,65,0,49.94,4934,0,Santa Monica,0,0,NA,34.035849,-118.50350800000001,1,20.05,0,7,None,11509,0,1,1,0,67,1,0.0,3345.98,43.66,1263.05,0,0,90402
3408,0,0,0,0,4,1,0,DSL,0,1,0,0,Month-to-month,0,Credit card (automatic),50.7,151.3,1,42,33,9.81,4930,1,Santa Monica,0,0,Cable,34.031529,-118.491156,0,52.728,0,0,None,23559,0,2,0,0,4,2,50.0,39.24,0.0,151.3,0,0,90403
3409,0,1,1,0,70,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,113.65,7714.65,0,77,25,35.39,6146,0,Santa Monica,1,0,Fiber Optic,34.026334000000006,-118.474222,1,113.65,0,7,None,19975,1,0,1,0,70,0,1929.0,2477.3,24.36,7714.65,0,0,90404
3410,1,0,0,0,3,1,0,DSL,0,0,1,0,Month-to-month,0,Credit card (automatic),53.4,188.7,1,23,90,47.68,2755,1,Santa Monica,0,1,Cable,34.005439,-118.477507,0,55.536,0,0,None,26099,0,1,0,1,3,2,170.0,143.04,0.0,188.7,1,0,90405
3411,1,1,1,0,53,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.9,5549.4,1,69,7,7.94,5884,1,Torrance,0,1,Cable,33.833698999999996,-118.31438700000001,1,105.976,0,1,Offer B,40705,0,0,1,0,53,3,0.0,420.82,0.0,5549.4,0,1,90501
3412,1,0,1,1,2,1,0,DSL,1,1,0,0,Two year,0,Mailed check,59.5,130.5,0,49,53,42.55,5613,0,Torrance,0,1,Cable,33.833181,-118.29206200000002,1,59.5,4,8,Offer E,17058,1,0,1,0,2,1,69.0,85.1,0.0,130.5,0,0,90502
3413,0,0,1,1,29,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),87.8,2621.75,0,32,13,33.62,4780,0,Torrance,0,0,Fiber Optic,33.840399,-118.353714,1,87.8,2,1,None,41979,0,0,1,1,29,0,34.08,974.98,0.0,2621.75,0,1,90503
3414,0,0,0,0,47,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,41.9,1875.25,0,54,23,0.0,2540,0,Torrance,1,0,Fiber Optic,33.867257,-118.330794,0,41.9,0,0,Offer B,31678,1,0,0,0,47,0,0.0,0.0,0.0,1875.25,0,1,90504
3415,0,0,1,1,68,1,1,Fiber optic,0,0,1,0,One year,1,Electronic check,83.0,5685.8,1,42,6,44.24,4714,1,Torrance,0,0,DSL,33.807882,-118.34795700000001,1,86.32000000000002,0,1,None,34873,0,3,1,0,68,1,341.0,3008.32,0.0,5685.8,0,0,90505
3416,1,0,0,1,12,1,0,DSL,1,0,1,1,Month-to-month,1,Mailed check,69.85,837.5,0,41,29,27.07,5796,0,Whittier,0,1,Fiber Optic,34.007353,-118.03368300000001,0,69.85,1,0,Offer D,32050,0,0,0,1,12,0,243.0,324.8400000000001,0.0,837.5,0,0,90601
3417,0,0,1,1,8,1,0,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),56.3,401.5,0,24,59,31.86,3135,0,Whittier,0,0,Fiber Optic,33.972119,-118.02018799999999,1,56.3,1,10,None,26265,1,1,1,0,8,2,237.0,254.88,0.0,401.5,1,0,90602
3418,1,0,1,0,54,1,1,Fiber optic,1,1,1,1,Month-to-month,0,Electronic check,109.55,6118.95,0,35,29,49.9,6130,0,Whittier,1,1,Cable,33.945318,-117.992066,1,109.55,0,9,Offer B,19109,0,0,1,1,54,3,1774.0,2694.6,0.0,6118.95,0,0,90603
3419,1,0,1,1,69,1,0,Fiber optic,0,1,1,0,Two year,1,Mailed check,92.15,6480.9,0,56,56,20.32,5817,0,Whittier,0,1,Cable,33.929704,-118.01208000000001,1,92.15,3,2,Offer A,37887,1,0,1,0,69,2,3629.0,1402.08,0.0,6480.9,0,0,90604
3420,0,0,0,0,26,1,1,DSL,1,1,1,0,Month-to-month,1,Bank transfer (automatic),69.5,1800.05,0,54,10,25.4,3866,0,Whittier,0,0,Fiber Optic,33.960891,-118.03222199999999,0,69.5,0,0,Offer C,38181,0,0,0,0,26,1,0.0,660.4,0.0,1800.05,0,1,90605
3421,0,0,1,0,72,1,1,Fiber optic,1,1,0,0,Two year,1,Bank transfer (automatic),97.0,7104.2,0,27,42,38.79,6302,0,Whittier,1,0,Fiber Optic,33.976678,-118.065875,1,97.0,0,1,Offer A,32148,1,1,1,0,72,1,298.38,2792.88,0.0,7104.2,1,1,90606
3422,0,0,0,0,70,0,No phone service,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),58.35,4214.25,0,54,13,0.0,4093,0,Buena Park,1,0,Fiber Optic,33.845706,-118.012204,0,58.35,0,0,Offer A,44442,1,0,0,1,70,0,54.79,0.0,0.0,4214.25,0,1,90620
3423,1,0,0,1,1,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,50.6,50.6,1,47,14,11.86,3677,1,Buena Park,0,1,Cable,33.874224,-117.99336799999999,0,52.623999999999995,2,0,None,33528,0,0,0,0,1,0,0.0,11.86,0.0,50.6,0,0,90621
3424,1,0,0,0,10,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.5,863.1,1,55,2,12.78,4206,1,La Palma,0,1,Cable,33.850504,-118.039892,0,93.08,0,0,Offer D,15505,0,0,0,1,10,5,17.0,127.8,0.0,863.1,0,0,90623
3425,0,0,1,1,28,1,0,Fiber optic,0,0,0,0,One year,1,Bank transfer (automatic),70.4,1992.2,0,56,24,12.94,5195,0,Cypress,0,0,DSL,33.818477,-118.038307,1,70.4,2,6,Offer C,47344,0,0,1,0,28,0,478.0,362.32,0.0,1992.2,0,0,90630
3426,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.8,69.8,1,50,28,22.86,4154,1,La Habra,0,1,DSL,33.940619,-117.9513,0,72.592,0,0,None,67354,0,2,0,0,1,3,0.0,22.86,0.0,69.8,0,1,90631
3427,0,0,1,0,21,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.3,1948.35,0,60,8,27.66,2058,0,La Mirada,0,0,Cable,33.902045,-118.00896100000001,1,94.3,0,6,Offer D,47568,0,0,1,1,21,0,156.0,580.86,0.0,1948.35,0,0,90638
3428,1,1,1,0,51,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Bank transfer (automatic),93.8,4750.95,1,80,33,22.14,4788,1,Montebello,1,1,Fiber Optic,34.015217,-118.10996200000001,1,97.552,0,1,Offer B,62425,0,1,1,0,51,1,1568.0,1129.14,0.0,4750.95,0,0,90640
3429,0,0,1,1,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.55,1007.9,0,49,0,30.31,4670,0,Norwalk,0,0,NA,33.905963,-118.08263000000001,1,19.55,1,10,Offer B,103214,0,0,1,0,53,0,0.0,1606.4299999999996,0.0,1007.9,0,0,90650
3430,1,0,0,1,53,1,0,Fiber optic,1,1,0,1,One year,0,Electronic check,95.95,5036.9,0,38,56,33.74,4523,0,Pico Rivera,1,1,Fiber Optic,33.989523999999996,-118.089299,0,95.95,3,0,Offer B,63288,0,0,0,1,53,0,2821.0,1788.22,0.0,5036.9,0,0,90660
3431,1,0,1,0,24,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.05,2391.8,1,44,25,34.62,4766,1,Santa Fe Springs,1,1,Cable,33.933565,-118.062611,1,105.09200000000001,0,1,None,16271,0,0,1,1,24,2,598.0,830.8799999999999,0.0,2391.8,0,0,90670
3432,0,0,1,0,70,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),94.8,6859.05,0,30,59,26.47,5072,0,Stanton,1,0,DSL,33.801869,-117.99506799999999,1,94.8,0,7,Offer A,29694,1,0,1,1,70,0,404.68,1852.9,0.0,6859.05,0,1,90680
3433,1,0,0,0,61,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,107.75,6521.9,0,30,71,42.4,5364,0,Artesia,1,1,Fiber Optic,33.867593,-118.08063700000001,0,107.75,0,0,Offer B,16398,0,0,0,1,61,4,0.0,2586.4,0.0,6521.9,0,1,90701
3434,0,0,0,0,11,1,0,DSL,1,0,0,0,One year,1,Mailed check,54.6,617.85,0,21,41,1.16,2573,0,Cerritos,0,0,DSL,33.8681,-118.067402,0,54.6,0,0,Offer D,51556,1,0,0,0,11,0,253.0,12.76,0.0,617.85,1,0,90703
3435,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),71.3,157.75,0,53,3,6.74,2274,0,Avalon,0,1,Cable,33.391181,-118.421305,0,71.3,0,0,Offer E,3699,0,0,0,0,2,0,0.0,13.48,0.0,157.75,0,1,90704
3436,1,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.5,516.3,0,29,0,3.58,4761,0,Bellflower,0,1,NA,33.887676,-118.12728899999999,0,19.5,0,0,Offer C,72893,0,0,0,0,25,0,0.0,89.5,0.0,516.3,1,0,90706
3437,0,0,0,0,41,1,1,DSL,0,1,0,0,One year,1,Credit card (automatic),56.3,2364,0,40,8,36.47,2994,0,Harbor City,0,0,Cable,33.798266,-118.30023700000001,0,56.3,0,0,Offer B,24660,0,0,0,0,41,0,0.0,1495.27,0.0,2364.0,0,1,90710
3438,1,0,1,0,18,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.7,1687.95,1,53,22,31.49,2206,1,Lakewood,0,1,Fiber Optic,33.840524,-118.148403,1,98.488,0,1,Offer D,30173,0,0,1,1,18,3,0.0,566.8199999999998,0.0,1687.95,0,1,90712
3439,1,1,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),104.15,7689.95,1,66,2,6.03,5925,1,Lakewood,1,1,DSL,33.847755,-118.112532,1,108.31600000000002,0,0,None,27563,0,0,0,0,72,2,154.0,434.16,0.0,7689.95,0,0,90713
3440,0,0,1,1,71,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),90.55,6239.05,0,43,20,41.71,6009,0,Lakewood,1,0,DSL,33.841027000000004,-118.078097,1,90.55,3,10,Offer A,20890,1,0,1,1,71,2,124.78,2961.41,0.0,6239.05,0,1,90715
3441,0,0,1,1,34,1,0,DSL,1,1,0,0,One year,1,Mailed check,60.8,2042.05,0,34,16,49.58,4522,0,Hawaiian Gardens,1,0,Fiber Optic,33.830431,-118.07407099999999,1,60.8,1,7,Offer C,14852,0,0,1,0,34,1,0.0,1685.72,0.0,2042.05,0,1,90716
3442,1,0,0,0,29,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),98.8,2807.1,0,62,19,48.2,4580,0,Lomita,1,1,DSL,33.794209,-118.31735400000001,0,98.8,0,0,Offer C,21065,1,0,0,1,29,0,0.0,1397.8000000000004,0.0,2807.1,0,1,90717
3443,1,1,1,0,40,1,0,Fiber optic,1,1,1,0,One year,1,Credit card (automatic),98.15,4116.8,0,68,18,15.15,4332,0,Los Alamitos,1,1,Cable,33.794990000000006,-118.065591,1,98.15,0,2,None,21343,1,0,1,0,40,1,741.0,606.0,27.89,4116.8,0,0,90720
3444,1,0,1,0,36,0,No phone service,DSL,1,0,0,0,One year,0,Mailed check,35.35,1317.95,0,37,23,0.0,3314,0,Paramount,1,1,Cable,33.897121999999996,-118.164432,1,35.35,0,7,Offer C,55306,0,0,1,0,36,0,303.0,0.0,0.0,1317.95,0,0,90723
3445,0,0,1,0,46,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,103.15,4594.65,0,41,29,33.22,3517,0,San Pedro,0,0,Fiber Optic,33.736387,-118.28436299999998,1,103.15,0,3,Offer B,58639,1,0,1,1,46,3,1332.0,1528.12,0.0,4594.65,0,0,90731
3446,0,0,0,0,58,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,107.75,6332.75,0,51,19,46.7,5121,0,San Pedro,1,0,Fiber Optic,33.744119,-118.31448,0,107.75,0,0,Offer B,21279,0,0,0,1,58,1,0.0,2708.600000000001,0.0,6332.75,0,1,90732
3447,1,0,0,0,39,1,1,Fiber optic,0,1,0,0,One year,0,Credit card (automatic),81.4,3213.75,0,54,12,36.93,4104,0,Seal Beach,0,1,Fiber Optic,33.75462,-118.071128,0,81.4,0,0,Offer C,24180,0,0,0,0,39,0,0.0,1440.27,0.0,3213.75,0,1,90740
3448,1,0,1,1,4,1,0,DSL,0,0,0,1,Month-to-month,0,Credit card (automatic),61.45,229.55,1,44,23,27.24,2131,1,Sunset Beach,0,1,Fiber Optic,33.719221000000005,-118.073596,1,63.90800000000001,1,4,None,1107,1,0,1,1,4,1,53.0,108.96,0.0,229.55,0,0,90742
3449,0,0,1,1,52,1,1,Fiber optic,0,1,1,0,One year,1,Credit card (automatic),95.7,4976.15,0,53,20,8.16,4415,0,Surfside,1,0,Fiber Optic,33.728273,-118.08530400000001,1,95.7,3,8,Offer B,174,0,0,1,0,52,0,995.0,424.32,0.0,4976.15,0,0,90743
3450,1,1,1,0,70,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,104.8,7308.95,0,66,28,39.49,5291,0,Wilmington,1,1,Cable,33.782068,-118.26226299999999,1,104.8,0,3,None,53323,0,0,1,0,70,0,2047.0,2764.3,6.11,7308.95,0,0,90744
3451,1,1,1,0,65,1,0,Fiber optic,0,0,0,0,One year,1,Bank transfer (automatic),70.95,4555.2,0,76,20,28.68,4871,0,Carson,0,1,Fiber Optic,33.822295000000004,-118.26411,1,70.95,0,6,None,55486,0,0,1,0,65,1,0.0,1864.2,7.43,4555.2,0,1,90745
3452,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.95,44.95,0,61,13,13.63,3256,0,Carson,0,1,DSL,33.859171,-118.25227199999999,0,44.95,0,0,Offer E,25566,0,0,0,0,1,0,0.0,13.63,0.0,44.95,0,0,90746
3453,0,0,1,0,70,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,97.65,6982.5,0,21,26,16.66,4252,0,Long Beach,1,0,DSL,33.752524,-118.21073700000001,1,97.65,0,9,Offer A,38427,0,0,1,1,70,1,0.0,1166.2,0.0,6982.5,1,1,90802
3454,0,1,1,1,29,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Mailed check,35.65,1025.15,0,67,20,0.0,4107,0,Long Beach,1,0,Fiber Optic,33.760458,-118.129725,1,35.65,1,8,None,31352,0,1,1,0,29,2,20.5,0.0,25.07,1025.15,0,1,90803
3455,1,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.55,90.55,1,20,53,7.15,3898,1,Long Beach,0,1,Cable,33.783046999999996,-118.1486,0,94.17200000000001,0,0,Offer E,43467,0,1,0,1,1,5,0.0,7.15,0.0,90.55,1,0,90804
3456,0,0,0,0,67,1,1,DSL,1,0,1,1,Two year,1,Mailed check,85.25,5714.2,0,21,41,8.71,6322,0,Long Beach,1,0,Fiber Optic,33.864622,-118.179626,0,85.25,0,0,Offer A,91664,1,0,0,1,67,4,234.28,583.57,1.31,5714.2,1,1,90805
3457,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.5,19.5,0,57,0,33.02,5279,0,Long Beach,0,0,NA,33.802664,-118.179971,0,19.5,0,0,Offer E,49647,0,0,0,0,1,0,0.0,33.02,0.0,19.5,0,0,90806
3458,0,0,0,0,26,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),88.8,2274.35,1,58,24,38.09,4910,1,Long Beach,0,0,DSL,33.830099,-118.182239,0,92.352,0,0,None,31556,0,2,0,1,26,4,546.0,990.34,0.0,2274.35,0,0,90807
3459,0,0,1,1,30,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,25.1,789.55,0,39,0,47.21,5851,0,Long Beach,0,0,NA,33.823943,-118.11133500000001,1,25.1,2,6,Offer C,37417,0,0,1,0,30,0,0.0,1416.3,15.41,789.55,0,0,90808
3460,0,0,1,0,48,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),100.05,4834,0,58,2,1.02,3468,0,Long Beach,1,0,Fiber Optic,33.819814,-118.222416,1,100.05,0,3,Offer B,35656,1,0,1,1,48,3,0.0,48.96,37.45,4834.0,0,1,90810
3461,0,0,1,1,55,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,55.7,3131.8,0,49,14,36.41,4149,0,Long Beach,0,0,Cable,33.781086,-118.199049,1,55.7,2,9,Offer B,63136,0,0,1,0,55,1,0.0,2002.55,34.16,3131.8,0,1,90813
3462,1,0,0,0,7,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Mailed check,85.2,602.55,1,23,29,18.83,3905,1,Long Beach,0,1,Cable,33.771612,-118.14386599999999,0,88.60799999999999,0,0,Offer E,19034,0,0,0,1,7,3,175.0,131.81,0.0,602.55,1,0,90814
3463,1,0,0,0,37,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Electronic check,91.15,3369.25,0,29,69,12.69,3194,0,Long Beach,0,1,DSL,33.797638,-118.11662,0,91.15,0,0,Offer C,38902,0,1,0,0,37,3,0.0,469.53,17.5,3369.25,1,1,90815
3464,0,0,1,0,31,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),83.85,2674.15,0,64,9,12.03,4283,0,Long Beach,0,0,Fiber Optic,33.778436,-118.118648,1,83.85,0,1,Offer C,425,0,0,1,1,31,3,0.0,372.93,11.37,2674.15,0,1,90822
3465,1,0,0,0,4,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.9,199.75,0,46,20,33.93,3200,0,Altadena,0,1,Fiber Optic,34.196837,-118.14223600000001,0,45.9,0,0,Offer E,36243,0,2,0,0,4,1,0.0,135.72,0.0,199.75,0,1,91001
3466,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.1,1790.8,0,49,0,27.93,4185,0,Arcadia,0,1,NA,34.137319,-118.02983700000001,1,25.1,2,7,Offer A,30028,0,0,1,0,72,1,0.0,2010.96,46.81,1790.8,0,0,91006
3467,1,1,0,0,5,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,91.4,449.75,1,79,12,4.59,2834,1,Arcadia,0,1,Fiber Optic,34.128284,-118.04773200000001,0,95.056,0,0,None,30933,0,2,0,0,5,3,0.0,22.95,0.0,449.75,0,1,91007
3468,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.7,19.7,0,37,0,34.28,2004,0,Duarte,0,1,NA,34.145695,-117.95982,1,19.7,3,2,None,27414,0,0,1,0,1,1,0.0,34.28,0.0,19.7,0,0,91010
3469,0,1,0,0,15,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,91.5,1400.3,0,80,16,39.57,4173,0,La Canada Flintridge,0,0,Cable,34.234912,-118.153729,0,91.5,0,0,None,20200,0,0,0,0,15,0,0.0,593.55,48.66,1400.3,0,1,91011
3470,1,0,1,1,8,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),51.3,411.6,0,47,20,10.36,2545,0,Monrovia,0,1,Fiber Optic,34.1528,-118.000482,1,51.3,1,7,None,41067,0,0,1,0,8,2,82.0,82.88,15.02,411.6,0,0,91016
3471,0,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,21.1,741,0,61,0,23.77,5707,0,Montrose,0,0,NA,34.2112,-118.230625,0,21.1,0,0,Offer C,7527,0,0,0,0,35,0,0.0,831.9499999999998,14.23,741.0,0,0,91020
3472,0,1,0,0,56,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,104.75,5841.35,0,67,7,27.64,5128,0,Sierra Madre,1,0,DSL,34.168686,-118.057505,0,104.75,0,0,None,10558,0,0,0,0,56,3,409.0,1547.84,36.52,5841.35,0,0,91024
3473,1,0,1,0,42,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),106.15,4512.7,1,54,23,2.41,2265,1,South Pasadena,1,1,Cable,34.110444,-118.156957,1,110.39600000000002,0,1,None,23984,1,3,1,1,42,1,1038.0,101.22,0.0,4512.7,0,0,91030
3474,1,1,1,1,65,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,85.75,5688.45,0,78,23,9.68,4978,0,Sunland,0,1,Fiber Optic,34.282703999999995,-118.312929,1,85.75,1,10,None,18752,0,0,1,0,65,2,0.0,629.1999999999998,38.09,5688.45,0,1,91040
3475,0,0,1,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.3,31.9,0,57,0,35.42,2843,0,Tujunga,0,0,NA,34.296574,-118.24483899999998,1,20.3,2,2,None,26753,0,0,1,0,2,1,0.0,70.84,0.0,31.9,0,0,91042
3476,1,1,1,0,65,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,100.75,6674.65,0,66,8,32.08,4368,0,Pasadena,0,1,Cable,34.146634999999996,-118.139225,1,100.75,0,6,None,16812,0,0,1,0,65,0,0.0,2085.2,0.0,6674.65,0,1,91101
3477,0,0,0,0,18,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.15,1345.75,0,43,13,11.36,5033,0,Pasadena,0,0,Cable,34.167465,-118.165327,0,74.15,0,0,Offer D,27891,0,0,0,0,18,0,0.0,204.48,0.0,1345.75,0,1,91103
3478,0,0,0,0,23,1,1,DSL,1,0,1,1,One year,1,Electronic check,78.55,1843.05,0,43,12,48.88,3127,0,Pasadena,1,0,DSL,34.165383,-118.123752,0,78.55,0,0,None,38460,0,0,0,1,23,0,221.0,1124.24,19.63,1843.05,0,0,91104
3479,0,0,0,0,4,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.3,196.95,1,36,22,39.9,3443,1,Pasadena,0,0,Fiber Optic,34.13946,-118.16664899999999,0,47.111999999999995,0,0,Offer E,10253,0,0,0,0,4,3,43.0,159.6,0.0,196.95,0,0,91105
3480,1,0,1,0,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.85,1433.8,0,30,0,3.51,4442,0,Pasadena,0,1,NA,34.139402000000004,-118.128658,1,19.85,0,9,Offer A,23742,0,0,1,0,70,2,0.0,245.7,45.47,1433.8,0,0,91106
3481,0,0,0,0,4,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,50.7,214.55,0,24,51,16.25,4288,0,Pasadena,0,0,Fiber Optic,34.159007,-118.08735300000001,0,50.7,0,0,None,32369,0,0,0,0,4,1,0.0,65.0,39.92,214.55,1,1,91107
3482,1,0,0,0,19,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),45.0,865.85,0,53,5,29.52,4519,0,San Marino,0,1,DSL,34.122671000000004,-118.11291100000001,0,45.0,0,0,None,13158,0,0,0,0,19,0,43.0,560.88,22.55,865.85,0,0,91108
3483,0,0,0,0,18,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,77.8,1358.6,0,61,26,19.93,4228,0,Glendale,1,0,DSL,34.17051,-118.28946299999998,0,77.8,0,0,None,23981,0,0,0,0,18,2,0.0,358.74,29.76,1358.6,0,1,91201
3484,0,1,1,0,38,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,83.45,3147.15,0,76,15,3.42,2768,0,Glendale,0,0,Fiber Optic,34.167926,-118.26753899999999,1,83.45,0,0,None,21990,0,1,0,0,38,1,472.0,129.96,24.98,3147.15,0,0,91202
3485,1,0,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),73.25,131.05,1,37,16,2.96,2919,1,Glendale,0,1,Cable,34.153338,-118.262974,0,76.18,0,0,None,14493,0,0,0,0,2,1,21.0,5.92,0.0,131.05,0,0,91203
3486,1,0,0,0,47,1,1,Fiber optic,1,1,1,0,One year,0,Bank transfer (automatic),94.8,4535.85,0,51,20,40.25,5022,0,Glendale,0,1,Fiber Optic,34.136306,-118.26036,0,94.8,0,0,Offer B,17015,0,0,0,0,47,1,90.72,1891.75,3.34,4535.85,0,1,91204
3487,0,0,1,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.1,1078.75,0,22,0,2.44,4529,0,Glendale,0,0,NA,34.13658,-118.24583899999999,1,20.1,1,10,None,41390,0,0,1,0,52,3,0.0,126.88,17.05,1078.75,1,0,91205
3488,1,0,0,0,9,1,1,DSL,0,0,0,1,Month-to-month,0,Mailed check,59.9,542.4,0,46,10,10.69,5414,0,Glendale,0,1,Fiber Optic,34.162515,-118.203869,0,59.9,0,0,None,31297,0,0,0,1,9,0,0.0,96.21,38.33,542.4,0,1,91206
3489,0,0,1,0,26,1,1,DSL,1,1,1,1,One year,1,Credit card (automatic),90.1,2312.55,0,46,19,25.63,2068,0,Glendale,1,0,Cable,34.182378,-118.262922,1,90.1,0,1,Offer C,9864,1,0,1,1,26,0,0.0,666.38,47.79,2312.55,0,1,91207
3490,1,0,1,1,8,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,51.05,415.05,1,47,22,3.85,3758,1,Glendale,1,1,DSL,34.195386,-118.23850800000001,1,53.092,1,1,Offer E,16910,0,3,1,0,8,2,0.0,30.8,0.0,415.05,0,1,91208
3491,1,0,1,0,44,1,0,DSL,0,1,1,0,One year,1,Electronic check,70.95,3250.45,0,19,48,29.61,3678,0,La Crescenta,1,1,Fiber Optic,34.239636,-118.245259,1,70.95,0,1,None,29110,1,0,1,0,44,0,0.0,1302.84,24.92,3250.45,1,1,91214
3492,0,0,0,0,3,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Mailed check,29.2,98.5,0,34,22,0.0,4699,0,Agoura Hills,0,0,DSL,34.129058,-118.75978799999999,0,29.2,0,0,None,25303,0,0,0,0,3,3,22.0,0.0,0.0,98.5,0,0,91301
3493,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),46.6,87.9,0,45,12,1.87,5096,0,Calabasas,0,1,Fiber Optic,34.130860999999996,-118.68346000000001,0,46.6,0,0,None,23661,0,0,0,0,2,0,11.0,3.74,0.0,87.9,0,0,91302
3494,0,0,1,1,9,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),85.35,754.65,1,63,6,14.21,2445,1,Canoga Park,0,0,DSL,34.19829,-118.602203,1,88.764,0,1,Offer E,23519,0,2,1,0,9,5,45.0,127.89,0.0,754.65,0,0,91303
3495,1,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.35,75.35,1,80,20,28.49,4403,1,Canoga Park,0,1,Cable,34.224377000000004,-118.63265600000001,0,78.36399999999998,0,0,None,49242,0,0,0,0,1,4,0.0,28.49,0.0,75.35,0,0,91304
3496,1,0,0,0,25,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Bank transfer (automatic),74.3,1952.25,0,53,26,17.3,4815,0,Winnetka,0,1,DSL,34.209532,-118.57756299999998,0,74.3,0,0,Offer C,43857,0,0,0,0,25,0,508.0,432.5,40.54,1952.25,0,0,91306
3497,0,1,1,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.3,153.8,0,79,2,32.62,2901,0,West Hills,0,0,DSL,34.199787,-118.68493000000001,1,69.3,0,1,Offer E,23637,0,0,1,0,2,0,3.0,65.24,0.0,153.8,0,0,91307
3498,1,0,0,0,43,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,75.2,3198.6,1,63,12,34.0,4673,1,Chatsworth,0,1,Cable,34.294142,-118.60388300000001,0,78.20800000000001,0,0,None,35325,0,2,0,0,43,2,384.0,1462.0,0.0,3198.6,0,0,91311
3499,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.9,20.9,1,54,0,15.51,5527,1,Encino,0,0,NA,34.150354,-118.51829199999999,0,20.9,0,0,Offer E,27614,0,0,0,0,1,0,0.0,15.51,0.0,20.9,0,0,91316
3500,0,0,1,0,58,1,1,Fiber optic,0,1,0,1,One year,1,Electronic check,94.3,5610.15,0,49,26,21.38,6166,0,Newbury Park,1,0,DSL,34.172071,-118.946262,1,94.3,0,1,None,37779,0,0,1,1,58,1,1459.0,1240.04,5.55,5610.15,0,0,91320
3501,0,0,1,1,59,1,1,DSL,1,0,1,0,Two year,1,Mailed check,76.45,4519.5,0,33,15,13.27,5978,0,Newhall,1,0,Fiber Optic,34.370378,-118.50411799999999,1,76.45,1,0,None,30742,1,0,0,0,59,1,0.0,782.93,30.22,4519.5,0,1,91321
3502,1,0,0,0,44,0,No phone service,DSL,1,0,1,1,One year,1,Electronic check,54.0,2440.25,0,55,17,0.0,4256,0,Northridge,1,1,DSL,34.238208,-118.55028999999999,0,54.0,0,0,None,25751,0,0,0,1,44,0,415.0,0.0,5.47,2440.25,0,0,91324
3503,1,0,0,0,66,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,104.25,6860.6,0,43,6,33.02,4915,0,Northridge,0,1,Fiber Optic,34.236683,-118.51758799999999,0,104.25,0,0,Offer A,32307,1,0,0,1,66,0,412.0,2179.32,44.0,6860.6,0,0,91325
3504,1,0,1,1,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.95,1377.7,0,45,0,35.89,4165,0,Porter Ranch,0,1,NA,34.281911,-118.55621799999999,1,19.95,3,1,Offer A,28067,0,0,1,0,68,0,0.0,2440.52,28.98,1377.7,0,0,91326
3505,1,0,0,0,9,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.95,190.25,0,61,7,0.0,5473,0,Pacoima,0,1,Fiber Optic,34.255441999999995,-118.421314,0,24.95,0,0,None,97318,0,0,0,0,9,0,13.0,0.0,0.0,190.25,0,0,91331
3506,1,0,0,0,19,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,84.75,1651.95,0,29,41,11.42,5157,0,Reseda,1,1,DSL,34.200175,-118.540958,0,84.75,0,0,None,68018,0,0,0,0,19,2,677.0,216.98,49.38,1651.95,1,0,91335
3507,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.75,78.3,0,20,0,41.94,4987,0,San Fernando,0,1,NA,34.286131,-118.435969,0,19.75,0,0,None,33389,0,0,0,0,4,0,0.0,167.76,0.0,78.3,1,0,91340
3508,0,0,0,0,70,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),113.65,7939.25,0,28,30,17.32,6424,0,Sylmar,1,0,DSL,34.321621,-118.399841,0,113.65,0,0,Offer A,81986,1,0,0,1,70,2,238.18,1212.4,0.0,7939.25,1,1,91342
3509,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.9,44.9,0,44,13,15.76,2451,0,North Hills,0,1,Fiber Optic,34.238802,-118.48229599999999,0,44.9,0,0,Offer E,57017,0,0,0,0,1,0,0.0,15.76,0.0,44.9,0,0,91343
3510,0,0,0,0,8,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.25,576.7,0,51,3,18.82,2332,0,Granada Hills,0,0,Fiber Optic,34.291273,-118.505104,0,75.25,0,0,None,48867,0,0,0,0,8,1,0.0,150.56,0.0,576.7,0,1,91344
3511,1,0,0,0,53,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.6,1279,0,24,0,34.16,4610,0,Mission Hills,0,1,NA,34.266389000000004,-118.459744,0,24.6,0,0,None,17112,0,0,0,0,53,2,0.0,1810.48,37.68,1279.0,1,0,91345
3512,1,1,0,0,51,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),25.0,1260.7,0,67,0,3.11,5896,0,Santa Clarita,0,1,NA,34.502432,-118.41458999999999,0,25.0,0,0,None,40077,0,0,0,0,51,0,0.0,158.61,0.0,1260.7,0,0,91350
3513,1,0,1,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.95,267.35,0,33,0,15.73,4075,0,Canyon Country,0,1,NA,34.422519,-118.420717,1,20.95,2,1,None,59259,0,0,1,0,11,0,0.0,173.03,18.17,267.35,0,0,91351
3514,1,0,1,1,60,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,110.6,6586.85,0,48,76,40.36,5756,0,Sun Valley,1,1,Fiber Optic,34.231053,-118.338307,1,110.6,3,1,None,46639,1,2,1,1,60,2,5006.0,2421.6,36.38,6586.85,0,0,91352
3515,1,0,0,0,17,1,0,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),55.5,934.15,0,64,14,33.68,3190,0,Valencia,0,1,Fiber Optic,34.457005,-118.57372600000001,0,55.5,0,0,None,17846,0,0,0,0,17,2,131.0,572.56,0.0,934.15,0,0,91354
3516,1,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,43.3,123.65,1,23,45,48.84,4849,1,Valencia,0,1,Cable,34.43987,-118.644609,0,45.032,0,0,Offer E,24977,0,2,0,1,3,6,56.0,146.52,0.0,123.65,1,0,91355
3517,1,0,1,0,70,1,0,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),109.5,7534.65,1,38,29,39.63,6136,1,Tarzana,1,1,Fiber Optic,34.157137,-118.548511,1,113.88,0,1,None,27424,1,0,1,1,70,1,2185.0,2774.100000000001,0.0,7534.65,0,0,91356
3518,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.45,19.45,0,34,0,29.15,2133,0,Thousand Oaks,0,1,NA,34.214054,-118.88108999999999,0,19.45,0,0,Offer E,42526,0,0,0,0,1,0,0.0,29.15,0.0,19.45,0,0,91360
3519,1,1,0,0,43,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.85,3645.6,0,74,7,8.81,4556,0,Westlake Village,0,1,Fiber Optic,34.130992,-118.894673,0,84.85,0,0,None,18735,0,0,0,0,43,0,255.0,378.83,0.0,3645.6,0,0,91361
3520,0,0,1,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.6,314.45,0,48,0,46.86,4298,0,Thousand Oaks,0,0,NA,34.191842,-118.822796,1,19.6,0,1,None,33057,0,1,1,0,16,1,0.0,749.76,26.83,314.45,0,0,91362
3521,0,0,1,1,57,1,0,DSL,1,1,0,0,One year,0,Electronic check,53.45,3053,0,33,11,17.01,5660,0,Woodland Hills,0,0,DSL,34.153733,-118.59340800000001,1,53.45,2,1,None,25988,0,0,1,0,57,1,33.58,969.57,0.0,3053.0,0,1,91364
3522,1,0,1,1,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.8,677.05,0,31,0,43.68,5137,0,Woodland Hills,0,1,NA,34.178067999999996,-118.61571399999998,1,19.8,1,1,None,36123,0,0,1,0,37,0,0.0,1616.16,29.21,677.05,0,0,91367
3523,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),112.1,7965.95,0,56,18,4.56,4272,0,Oak Park,1,0,DSL,34.19225,-118.77687399999999,1,112.1,0,1,None,14814,1,0,1,1,72,2,1434.0,328.32,18.88,7965.95,0,0,91377
3524,0,1,0,0,11,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),84.8,906.85,1,78,6,4.1,5118,1,Stevenson Ranch,0,0,Fiber Optic,34.364153,-118.615583,0,88.19200000000001,0,0,None,9937,0,0,0,0,11,0,0.0,45.1,0.0,906.85,0,1,91381
3525,0,1,1,0,50,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,95.05,4888.7,1,67,4,31.56,5863,1,Castaic,1,0,Fiber Optic,34.506627,-118.699048,1,98.852,0,1,Offer B,22177,0,2,1,0,50,1,0.0,1578.0,0.0,4888.7,0,1,91384
3526,1,1,0,0,5,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,50.35,237.25,1,73,31,18.69,4618,1,Van Nuys,1,1,DSL,34.178483,-118.43179099999999,0,52.364,0,0,None,40376,0,1,0,0,5,3,74.0,93.45,0.0,237.25,0,0,91401
3527,1,0,1,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.6,74.6,1,63,3,44.73,5861,1,Fallbrook,0,1,Fiber Optic,33.362575,-117.299644,1,77.584,0,1,Offer E,42239,0,0,1,0,1,2,0.0,44.73,0.0,74.6,0,0,92028
3528,1,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.7,342.4,1,35,0,5.74,3438,1,Sherman Oaks,0,1,NA,34.147149,-118.463365,0,19.7,0,0,Offer D,22085,0,0,0,0,16,0,0.0,91.84,0.0,342.4,0,0,91403
3529,1,1,1,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.2,140.1,0,69,14,7.29,3170,0,Van Nuys,1,1,Cable,34.202494,-118.448048,1,74.2,0,1,Offer E,51348,0,0,1,0,2,0,0.0,14.58,0.0,140.1,0,1,91405
3530,0,0,0,0,17,1,1,DSL,0,0,1,0,Month-to-month,1,Mailed check,69.0,1108,0,53,14,5.49,4439,0,Van Nuys,1,0,Fiber Optic,34.195685,-118.490752,0,69.0,0,0,None,50047,1,0,0,0,17,2,155.0,93.33,33.67,1108.0,0,0,91406
3531,0,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.35,295.55,0,63,0,40.95,2017,0,Van Nuys,0,0,NA,34.178470000000004,-118.45947199999999,0,19.35,0,0,None,23646,0,0,0,0,16,0,0.0,655.2,0.0,295.55,0,0,91411
3532,0,0,0,0,15,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,59.45,892.65,1,25,53,36.34,5129,1,Sherman Oaks,1,0,Cable,34.146957,-118.432138,0,61.828,0,0,Offer D,29387,0,0,0,1,15,0,473.0,545.1,0.0,892.65,1,0,91423
3533,0,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.8,198.25,0,57,0,2.84,5270,0,Encino,0,0,NA,34.152875,-118.486056,0,19.8,0,0,None,13129,0,0,0,0,10,0,0.0,28.4,0.0,198.25,0,0,91436
3534,0,0,0,1,46,1,0,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),105.2,4822.85,1,23,78,43.04,3322,1,Burbank,0,0,DSL,34.188339,-118.30094199999999,0,109.40799999999999,0,0,None,18112,1,0,0,1,46,2,0.0,1979.84,0.0,4822.85,1,1,91501
3535,1,0,1,1,64,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),109.2,6741.15,0,53,12,13.73,5543,0,Burbank,1,1,Fiber Optic,34.177267,-118.31003,1,109.2,1,1,None,11517,1,0,1,1,64,0,809.0,878.72,17.3,6741.15,0,0,91502
3536,0,0,0,0,1,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,79.15,79.15,0,33,23,18.0,2742,0,Burbank,0,0,Fiber Optic,34.213049,-118.317651,0,79.15,0,0,Offer E,25882,0,1,0,0,1,1,0.0,18.0,0.0,79.15,0,1,91504
3537,1,0,1,1,25,1,0,DSL,0,1,0,0,One year,0,Mailed check,53.65,1355.45,0,63,53,36.17,5854,0,Burbank,1,1,Fiber Optic,34.174215000000004,-118.345928,1,53.65,3,1,None,29245,0,0,1,0,25,1,718.0,904.25,0.0,1355.45,0,0,91505
3538,1,0,1,1,71,1,0,Fiber optic,1,1,1,0,Two year,0,Credit card (automatic),100.2,7209,0,22,27,33.69,5502,0,Burbank,1,1,DSL,34.169706,-118.323548,1,100.2,1,1,None,18539,1,0,1,0,71,0,0.0,2391.99,0.0,7209.0,1,1,91506
3539,1,0,0,0,8,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.15,438.4,1,59,6,35.53,3721,1,Los Angeles,0,1,DSL,34.099869,-118.326843,0,46.956,0,0,None,30568,0,0,0,0,8,3,26.0,284.24,0.0,438.4,0,0,90028
3540,0,0,1,1,72,1,0,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),108.65,7726.35,0,63,29,14.46,5730,0,North Hollywood,1,0,Cable,34.15136,-118.36478600000001,1,108.65,1,1,None,16996,1,0,1,1,72,0,0.0,1041.12,0.0,7726.35,0,1,91602
3541,0,0,1,0,49,0,No phone service,DSL,1,0,1,0,Month-to-month,0,Bank transfer (automatic),40.65,2070.75,0,57,11,0.0,5565,0,Studio City,0,0,Cable,34.139082,-118.39275,1,40.65,0,6,None,26157,0,0,1,0,49,1,0.0,0.0,0.0,2070.75,0,1,91604
3542,1,0,1,1,29,0,No phone service,DSL,1,1,0,1,One year,1,Credit card (automatic),55.35,1636.95,0,62,57,0.0,5138,0,North Hollywood,1,1,Fiber Optic,34.207295,-118.40002199999999,1,55.35,3,6,None,57146,1,0,1,1,29,0,933.0,0.0,0.0,1636.95,0,0,91605
3543,1,0,1,0,72,1,1,Fiber optic,1,1,0,1,Two year,0,Bank transfer (automatic),105.6,7581.5,0,59,5,6.15,5981,0,North Hollywood,1,1,Cable,34.187599,-118.387125,1,105.6,0,5,None,45358,1,1,1,1,72,3,0.0,442.8,0.0,7581.5,0,1,91606
3544,1,0,1,0,31,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Electronic check,93.8,3019.5,1,62,19,2.12,4115,1,Valley Village,1,1,DSL,34.165783000000005,-118.399795,1,97.552,0,1,None,27453,0,1,1,0,31,1,574.0,65.72,0.0,3019.5,0,0,91607
3545,0,0,0,0,50,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.7,4729.75,0,42,6,49.14,4164,0,Rancho Cucamonga,0,0,Cable,34.132275,-117.611478,0,95.7,0,0,None,39064,0,0,0,1,50,2,0.0,2457.0,0.0,4729.75,0,1,91701
3546,1,0,1,0,71,1,1,DSL,1,0,1,1,Two year,0,Electronic check,83.2,6126.1,0,47,12,35.09,5350,0,Azusa,1,1,Cable,34.174493,-117.87068000000001,1,83.2,0,6,None,57775,1,0,1,1,71,2,735.0,2491.390000000001,0.0,6126.1,0,0,91702
3547,1,1,1,0,70,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),90.05,6333.4,0,65,17,12.07,4666,0,Baldwin Park,1,1,Fiber Optic,34.098275,-117.967399,1,90.05,0,7,None,76890,1,0,1,1,70,0,1077.0,844.9,0.0,6333.4,0,0,91706
3548,1,0,0,0,71,1,1,Fiber optic,1,0,0,1,One year,0,Credit card (automatic),97.65,6687.85,0,47,5,16.57,5319,0,Chino Hills,0,1,Fiber Optic,33.942895,-117.72564399999999,0,97.65,0,0,None,66754,1,0,0,1,71,1,334.0,1176.47,0.0,6687.85,0,0,91709
3549,1,0,1,1,61,1,0,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),68.05,4158.25,0,23,59,42.31,4436,0,Chino,1,1,DSL,33.990646000000005,-117.663025,1,68.05,2,2,None,75319,1,0,1,0,61,1,0.0,2580.9100000000008,0.0,4158.25,1,1,91710
3550,1,0,0,0,32,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.2,3183.4,1,45,29,25.21,3606,1,Claremont,0,1,DSL,34.127621000000005,-117.717863,0,100.04799999999999,0,0,None,34716,1,0,0,1,32,4,923.0,806.72,0.0,3183.4,0,0,91711
3551,0,0,0,1,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.6,79.6,1,20,57,21.72,3108,1,Covina,0,0,Cable,34.097345000000004,-117.90673600000001,0,82.78399999999998,0,0,Offer E,33817,0,2,0,1,1,1,0.0,21.72,0.0,79.6,1,0,91722
3552,1,0,0,0,68,1,1,Fiber optic,1,1,0,1,Two year,1,Bank transfer (automatic),102.1,7149.35,0,40,7,49.42,5228,0,Covina,1,1,DSL,34.084747,-117.886844,0,102.1,0,0,None,17554,0,0,0,1,68,0,0.0,3360.56,0.0,7149.35,0,1,91723
3553,1,0,0,0,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),23.4,1429.65,0,43,0,48.93,5822,0,Covina,0,1,NA,34.081109999999995,-117.853935,0,23.4,0,0,None,25068,0,0,0,0,62,1,0.0,3033.66,0.0,1429.65,0,0,91724
3554,0,0,0,1,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.05,472.65,0,48,13,28.5,4668,0,Rancho Cucamonga,0,0,Fiber Optic,34.100970000000004,-117.57882,0,71.05,1,0,Offer E,51970,0,0,0,0,7,2,0.0,199.5,0.0,472.65,0,1,91730
3555,1,0,0,0,20,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.25,1734.5,1,49,28,1.36,2414,1,El Monte,0,1,Cable,34.079934,-118.046695,0,88.66,0,0,Offer D,30211,0,1,0,0,20,3,486.0,27.200000000000006,0.0,1734.5,0,0,91731
3556,1,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.45,113.5,0,53,0,1.57,3461,0,El Monte,0,1,NA,34.074492,-118.01462,1,19.45,3,10,Offer E,62660,0,0,1,0,6,1,0.0,9.42,0.0,113.5,0,0,91732
3557,0,1,0,0,33,0,No phone service,DSL,1,1,1,1,Month-to-month,1,Bank transfer (automatic),59.45,1884.65,0,80,16,0.0,3116,0,South El Monte,1,0,DSL,34.04622,-118.053753,0,59.45,0,0,None,45645,0,0,0,0,33,2,302.0,0.0,0.0,1884.65,0,0,91733
3558,1,0,1,1,28,1,1,Fiber optic,0,0,1,1,One year,0,Bank transfer (automatic),92.2,2568.15,0,37,30,13.19,5116,0,Rancho Cucamonga,0,1,DSL,34.245289,-117.642503,1,92.2,3,1,None,23079,0,0,1,1,28,0,77.04,369.32,0.0,2568.15,0,1,91737
3559,1,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.85,470,0,27,0,47.65,2176,0,Rancho Cucamonga,0,1,NA,34.133809,-117.523724,0,19.85,0,0,None,12937,0,0,0,0,27,2,0.0,1286.55,0.0,470.0,1,0,91739
3560,1,0,0,0,7,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,43.9,278.4,0,41,6,30.04,3565,0,Glendora,0,1,Fiber Optic,34.119363,-117.85505900000001,0,43.9,0,0,Offer E,25135,0,0,0,0,7,1,0.0,210.28,0.0,278.4,0,1,91740
3561,1,0,0,0,26,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,80.5,2088.8,1,34,24,24.16,2729,1,Glendora,0,1,Cable,34.14649,-117.84981499999999,0,83.72,0,0,None,24973,1,0,0,0,26,3,501.0,628.16,0.0,2088.8,0,0,91741
3562,1,1,0,0,5,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.8,502.6,1,75,13,36.36,2960,1,North Hollywood,0,1,Cable,34.207295,-118.40002199999999,0,93.39200000000001,0,0,None,57146,0,0,0,0,5,0,6.53,181.8,0.0,502.6,0,1,91605
3563,1,1,0,0,30,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Credit card (automatic),90.5,2595.85,0,69,14,4.04,5983,0,Hacienda Heights,0,1,Fiber Optic,33.998471,-117.973758,0,90.5,0,0,None,53686,0,0,0,0,30,0,363.0,121.2,0.0,2595.85,0,0,91745
3564,1,0,0,0,63,1,1,Fiber optic,0,1,0,1,One year,0,Credit card (automatic),90.45,5825.5,0,33,28,9.21,4616,0,La Puente,0,1,DSL,34.038983,-117.991372,0,90.45,0,0,None,30802,0,1,0,1,63,1,1631.0,580.23,0.0,5825.5,0,0,91746
3565,1,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,50.75,50.75,1,61,3,43.03,5355,1,Rowland Heights,0,1,DSL,33.976753,-117.89736699999999,0,52.78,0,0,Offer E,46342,0,1,0,0,1,2,0.0,43.03,0.0,50.75,0,0,91748
3566,0,0,0,1,53,1,1,DSL,0,1,1,1,One year,1,Electronic check,84.6,4449.75,0,55,18,14.54,4733,0,La Verne,1,0,Fiber Optic,34.144703,-117.770299,0,84.6,2,0,None,35530,1,0,0,1,53,2,0.0,770.62,0.0,4449.75,0,1,91750
3567,0,0,1,1,14,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),89.65,1208.35,1,57,3,7.62,2504,1,Mira Loma,0,0,DSL,33.999992,-117.535395,1,93.236,0,1,Offer D,18980,1,1,1,1,14,2,3.63,106.68,0.0,1208.35,0,1,91752
3568,0,0,0,0,21,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),99.15,1956.4,0,22,51,6.12,5324,0,Monterey Park,0,0,DSL,34.050321999999994,-118.14703700000001,0,99.15,0,0,Offer D,33280,1,0,0,1,21,2,998.0,128.52,0.0,1956.4,1,0,91754
3569,1,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.95,310.6,0,23,0,25.91,2221,0,Monterey Park,0,1,NA,34.049172,-118.115022,0,19.95,0,0,Offer D,26933,0,0,0,0,17,2,0.0,440.47,0.0,310.6,1,0,91755
3570,1,0,1,1,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.5,290.55,0,30,0,27.24,2856,0,Mt Baldy,0,1,NA,34.231318,-117.66203200000001,1,20.5,2,3,Offer D,47,0,0,1,0,16,0,0.0,435.84,0.0,290.55,0,0,91759
3571,0,0,0,0,35,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,62.1,2096.1,0,61,7,2.15,5315,0,Ontario,1,0,DSL,34.035602000000004,-117.591528,0,62.1,0,0,None,56280,0,0,0,1,35,2,147.0,75.25,0.0,2096.1,0,0,91761
3572,0,1,0,0,32,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.5,2665,0,74,12,48.62,3041,0,Ontario,0,0,Cable,34.057256,-117.667677,0,79.5,0,0,None,54254,0,2,0,0,32,1,31.98,1555.84,0.0,2665.0,0,1,91762
3573,0,0,1,1,28,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.55,543.8,0,27,0,15.85,3948,0,Montclair,0,0,NA,34.072121,-117.698319,1,19.55,3,9,None,34447,0,1,1,0,28,3,0.0,443.8,0.0,543.8,1,0,91763
3574,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.35,20.35,0,30,0,29.86,2183,0,Ontario,0,0,NA,34.074087,-117.60561799999999,0,20.35,0,0,Offer E,49474,0,2,0,0,1,1,0.0,29.86,0.0,20.35,0,0,91764
3575,1,0,0,0,59,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,51.7,3005.8,0,43,7,0.0,6107,0,Diamond Bar,0,1,Fiber Optic,33.992416,-117.807874,0,51.7,0,0,None,46532,1,0,0,1,59,2,210.0,0.0,0.0,3005.8,0,0,91765
3576,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),23.3,1623.15,0,26,0,18.14,4152,0,Pomona,0,0,NA,34.042286,-117.756106,1,23.3,2,6,None,69974,0,0,1,0,72,0,0.0,1306.08,0.0,1623.15,1,0,91766
3577,1,0,0,0,36,1,0,DSL,0,1,0,1,One year,1,Mailed check,65.4,2498.4,1,25,94,26.51,5220,1,Pomona,0,1,Cable,34.083086,-117.737997,0,68.016,0,0,None,46626,1,1,0,1,36,5,0.0,954.36,0.0,2498.4,1,1,91767
3578,0,0,0,0,40,1,0,DSL,1,1,1,0,Month-to-month,0,Mailed check,65.1,2586,0,32,26,11.56,3885,0,Pomona,0,0,DSL,34.067932,-117.785168,0,65.1,0,0,None,36057,0,0,0,0,40,2,0.0,462.4,0.0,2586.0,0,1,91768
3579,1,0,1,1,40,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,81.2,3292.3,0,55,56,3.52,5370,0,Rosemead,1,1,Fiber Optic,34.065108,-118.08279099999999,1,81.2,3,4,None,61623,0,0,1,0,40,1,0.0,140.8,0.0,3292.3,0,1,91770
3580,0,0,0,1,9,1,0,DSL,0,0,1,1,Month-to-month,1,Mailed check,72.9,651.4,1,50,12,35.49,3585,1,San Dimas,1,0,DSL,34.102119,-117.815532,0,75.816,2,0,None,33878,1,1,0,1,9,4,78.0,319.41,0.0,651.4,0,0,91773
3581,1,0,1,1,63,1,0,DSL,1,1,1,0,Two year,0,Credit card (automatic),74.5,4674.55,0,22,73,42.17,6382,0,San Gabriel,1,1,Cable,34.114771999999995,-118.089431,1,74.5,2,9,None,23444,1,0,1,0,63,1,0.0,2656.71,0.0,4674.55,1,1,91775
3582,0,0,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.5,232.35,0,48,5,26.86,2032,0,San Gabriel,0,0,DSL,34.089927,-118.09564499999999,0,80.5,0,0,None,38041,0,0,0,0,3,0,12.0,80.58,0.0,232.35,0,0,91776
3583,1,0,1,1,40,0,No phone service,DSL,0,1,1,1,One year,0,Mailed check,60.3,2448.5,0,19,26,0.0,3724,0,Temple City,1,1,Fiber Optic,34.101608,-118.055848,1,60.3,2,3,None,32718,1,0,1,1,40,0,0.0,0.0,0.0,2448.5,1,1,91780
3584,1,0,1,0,8,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,75.0,658.1,0,57,18,20.67,5413,0,Upland,0,1,DSL,34.141146,-117.65558300000001,1,75.0,0,8,Offer E,23331,0,0,1,0,8,2,118.0,165.36,0.0,658.1,0,0,91784
3585,1,1,1,0,34,1,0,Fiber optic,1,0,1,0,One year,0,Mailed check,90.15,3128.8,0,71,18,26.49,3202,0,Upland,0,1,Cable,34.105493,-117.66093400000001,1,90.15,0,7,None,48827,1,0,1,0,34,0,56.32,900.66,0.0,3128.8,0,1,91786
3586,1,0,0,0,5,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,40.0,223.45,1,25,65,0.0,3125,1,Walnut,1,1,Cable,34.018353999999995,-117.85491999999999,0,41.6,0,0,None,45118,1,3,0,1,5,2,0.0,0.0,0.0,223.45,1,1,91789
3587,1,1,0,0,9,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),99.45,919.4,1,67,16,10.66,2313,1,West Covina,0,1,DSL,34.066964,-117.93700700000001,0,103.428,0,0,None,44099,0,2,0,0,9,2,0.0,95.94,0.0,919.4,0,1,91790
3588,1,0,1,0,9,1,1,DSL,0,1,0,1,Month-to-month,1,Credit card (automatic),69.05,653.95,0,27,59,26.03,2907,0,West Covina,1,1,Cable,34.061634000000005,-117.893169,1,69.05,0,4,Offer E,30458,0,0,1,1,9,3,0.0,234.27,0.0,653.95,1,1,91791
3589,1,0,1,1,31,1,1,DSL,0,0,0,1,Month-to-month,0,Bank transfer (automatic),59.7,1825.5,0,21,59,30.67,2425,0,West Covina,0,1,Fiber Optic,34.024405,-117.89872199999999,1,59.7,1,6,None,31622,0,0,1,1,31,0,1077.0,950.77,0.0,1825.5,1,0,91792
3590,0,0,1,0,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.85,943.1,0,30,0,28.1,4358,0,Alhambra,0,0,NA,34.090925,-118.12816399999998,1,19.85,0,1,None,54382,0,0,1,0,50,1,0.0,1405.0,0.0,943.1,0,0,91801
3591,0,0,0,0,2,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,86.25,181.65,1,40,18,36.81,3529,1,Alhambra,0,0,Cable,34.074736,-118.145959,0,89.7,0,0,None,30635,1,0,0,0,2,0,33.0,73.62,0.0,181.65,0,0,91803
3592,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.65,45.65,1,43,24,36.99,4689,1,Alpine,0,0,Cable,32.827184,-116.70372900000001,0,47.476000000000006,0,0,None,16486,0,1,0,0,1,2,0.0,36.99,0.0,45.65,0,0,91901
3593,1,0,0,0,8,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.1,551.35,1,30,94,13.04,2899,1,Bonita,0,1,Cable,32.671170000000004,-117.00232,0,72.904,0,0,None,17389,0,0,0,0,8,1,518.0,104.32,0.0,551.35,0,0,91902
3594,0,0,0,0,9,0,No phone service,DSL,0,1,0,1,Month-to-month,0,Electronic check,40.75,359.4,0,45,21,0.0,2973,0,Boulevard,0,0,DSL,32.677096999999996,-116.30499099999999,0,40.75,0,0,Offer E,1509,0,0,0,1,9,0,75.0,0.0,0.0,359.4,0,0,91905
3595,0,1,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),70.2,115.95,1,75,31,9.55,2767,1,Campo,0,0,DSL,32.673483000000004,-116.47286299999999,0,73.00800000000002,0,0,None,3133,0,0,0,0,2,4,36.0,19.1,0.0,115.95,0,0,91906
3596,0,0,0,0,3,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,55.35,165.2,1,19,57,1.24,5787,1,Chula Vista,0,0,DSL,32.636792,-117.05498899999999,0,57.56399999999999,0,0,None,74025,0,1,0,1,3,3,94.0,3.72,0.0,165.2,1,0,91910
3597,1,0,1,0,25,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),95.7,2338.35,0,51,8,3.81,4535,0,Chula Vista,0,1,DSL,32.607964,-117.059459,1,95.7,0,7,None,71126,1,0,1,1,25,1,187.0,95.25,0.0,2338.35,0,0,91911
3598,1,1,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,46.3,46.3,0,71,21,11.51,2546,0,Chula Vista,0,1,Fiber Optic,32.64164,-116.985026,0,46.3,0,0,Offer E,12884,0,0,0,0,1,2,0.0,11.51,0.0,46.3,0,1,91913
3599,0,0,1,1,45,1,1,DSL,1,1,1,0,Month-to-month,0,Mailed check,81.3,3541.1,0,51,11,10.21,3111,0,Chula Vista,1,0,Fiber Optic,32.688506,-116.93863200000001,1,81.3,2,9,Offer B,2606,1,0,1,0,45,1,390.0,459.4500000000001,0.0,3541.1,0,0,91914
3600,1,1,1,1,51,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,84.2,4146.05,1,80,24,43.58,6245,1,Chula Vista,1,1,Cable,32.605012,-116.97595,1,87.56800000000001,0,2,Offer B,9278,0,0,1,0,51,1,0.0,2222.58,0.0,4146.05,0,1,91915
3601,0,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.0,1087.25,0,31,0,31.3,4277,0,Descanso,0,0,NA,32.912664,-116.63538700000001,1,20.0,1,4,Offer B,1587,0,0,1,0,55,2,0.0,1721.5,0.0,1087.25,0,0,91916
3602,0,0,0,0,38,1,1,DSL,1,1,0,0,Month-to-month,1,Bank transfer (automatic),66.15,2522.4,0,39,13,20.14,4933,0,Dulzura,1,0,DSL,32.622999,-116.687855,0,66.15,0,0,None,727,0,0,0,0,38,0,328.0,765.32,0.0,2522.4,0,0,91917
3603,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.85,81,1,34,18,19.52,3843,1,Guatay,0,1,DSL,32.857946000000005,-116.561917,0,47.68400000000001,0,0,None,796,0,0,0,0,2,1,15.0,39.04,0.0,81.0,0,0,91931
3604,1,0,1,1,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.6,717.3,0,40,0,24.16,3854,0,Imperial Beach,0,1,NA,32.579134,-117.119009,1,19.6,2,3,None,26662,0,0,1,0,38,1,0.0,918.08,0.0,717.3,0,0,91932
3605,1,0,0,0,34,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,49.8,1734.2,0,34,27,4.89,2711,0,Jacumba,0,1,DSL,32.649786999999996,-116.2237,0,49.8,0,0,None,699,0,0,0,0,34,0,468.0,166.26,0.0,1734.2,0,0,91934
3606,0,0,1,0,70,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,101.75,7069.3,0,19,26,19.88,5596,0,Jamul,1,0,Fiber Optic,32.695681,-116.79838600000001,1,101.75,0,0,None,8759,0,0,0,1,70,0,0.0,1391.6,0.0,7069.3,1,1,91935
3607,0,0,0,0,13,1,0,DSL,1,0,0,0,One year,0,Mailed check,55.15,742.9,0,20,59,46.68,3161,0,La Mesa,0,0,Fiber Optic,32.759327,-116.99726000000001,0,55.15,0,0,Offer D,44652,1,0,0,1,13,1,0.0,606.84,0.0,742.9,1,1,91941
3608,1,0,0,0,39,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.25,3017.65,1,64,6,36.17,4696,1,La Mesa,0,1,Cable,32.782501,-117.01611000000001,0,78.26,0,0,Offer C,24005,0,0,0,0,39,2,181.0,1410.63,0.0,3017.65,0,0,91942
3609,0,0,0,0,61,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,103.95,6423,0,21,30,15.44,4148,0,Lemon Grove,1,0,DSL,32.733564,-117.03371299999999,0,103.95,0,0,Offer B,24961,0,1,0,1,61,2,0.0,941.84,0.0,6423.0,1,1,91945
3610,0,0,0,0,12,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),100.15,1164.3,1,24,52,30.54,3682,1,Mount Laguna,1,0,Cable,32.830852,-116.444601,0,104.156,0,0,Offer D,81,0,0,0,1,12,5,605.0,366.48,0.0,1164.3,1,0,91948
3611,1,0,0,0,41,1,0,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),99.65,4220.35,0,29,59,21.64,2640,0,National City,0,1,Fiber Optic,32.67102,-117.095235,0,99.65,0,0,Offer B,62355,1,0,0,1,41,0,2490.0,887.24,0.0,4220.35,1,0,91950
3612,1,0,0,0,21,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.7,1558.7,0,28,42,28.54,2071,0,Pine Valley,0,1,Cable,32.800671,-116.48336299999998,0,73.7,0,0,Offer D,1604,0,0,0,1,21,0,0.0,599.34,0.0,1558.7,1,1,91962
3613,1,1,0,0,55,0,No phone service,DSL,0,0,1,1,One year,1,Bank transfer (automatic),50.05,2743.45,0,71,23,0.0,4932,0,Potrero,1,1,Fiber Optic,32.619465000000005,-116.59360500000001,0,50.05,0,0,None,905,0,0,0,0,55,2,631.0,0.0,0.0,2743.45,0,0,91963
3614,1,0,1,0,69,0,No phone service,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),60.25,4055.5,0,22,59,0.0,5717,0,Spring Valley,1,1,Fiber Optic,32.726627,-116.99460800000001,1,60.25,0,7,None,56100,1,0,1,1,69,1,0.0,0.0,0.0,4055.5,1,1,91977
3615,1,1,1,1,26,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,105.75,2710.25,1,72,20,1.26,3157,1,Spring Valley,1,1,DSL,32.730264,-116.95096299999999,1,109.98,0,0,Offer C,7863,0,4,0,1,26,3,542.0,32.76,0.0,2710.25,0,0,91978
3616,0,1,1,0,69,1,0,Fiber optic,1,1,0,1,One year,0,Credit card (automatic),87.3,6055.55,0,67,19,34.55,4148,0,Tecate,0,0,Cable,32.587557000000004,-116.636816,1,87.3,0,6,None,91,0,1,1,0,69,1,1151.0,2383.95,0.0,6055.55,0,0,91980
3617,0,1,1,0,18,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,48.35,810.7,1,70,13,0.0,2167,1,Bonsall,1,0,Cable,33.290907000000004,-117.202895,1,50.284000000000006,0,1,None,3849,0,3,1,1,18,1,105.0,0.0,0.0,810.7,0,0,92003
3618,1,0,1,1,47,1,1,DSL,0,1,0,0,Month-to-month,0,Electronic check,54.25,2538.2,0,28,26,39.25,2320,0,Borrego Springs,0,1,Fiber Optic,33.200369,-116.19231299999998,1,54.25,1,1,Offer B,2863,0,0,1,1,47,0,660.0,1844.75,0.0,2538.2,1,0,92004
3619,0,0,1,1,72,1,0,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),85.3,6129.2,0,46,21,36.13,4456,0,Cardiff By The Sea,1,0,Fiber Optic,33.015865999999995,-117.272254,1,85.3,1,0,None,10375,1,0,0,1,72,1,0.0,2601.36,0.0,6129.2,0,1,92007
3620,1,1,1,0,33,0,No phone service,DSL,0,1,1,0,Month-to-month,1,Electronic check,50.0,1750.85,0,80,4,0.0,5600,0,Carlsbad,1,1,DSL,33.148115999999995,-117.30604299999999,1,50.0,0,1,None,35582,1,0,1,0,33,0,70.0,0.0,0.0,1750.85,0,0,92008
3621,0,0,1,1,2,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,24.4,36.55,1,53,57,0.0,2635,1,Carlsbad,0,0,Cable,33.098017999999996,-117.25820300000001,1,25.376,3,0,None,43161,0,0,0,0,2,2,0.0,0.0,0.0,36.55,0,1,92009
3622,0,0,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),90.95,6652.45,0,20,47,45.66,5096,0,Del Mar,1,0,DSL,32.948262,-117.25608600000001,1,90.95,1,2,None,13945,1,0,1,1,72,1,3127.0,3287.5199999999995,0.0,6652.45,1,0,92014
3623,1,1,1,0,37,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),72.25,2575.45,0,75,7,23.54,4121,0,El Cajon,0,1,Fiber Optic,32.785165,-116.862648,1,72.25,0,8,None,40995,0,0,1,0,37,2,0.0,870.98,0.0,2575.45,0,1,92019
3624,0,1,1,1,62,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),96.1,6019.35,0,67,12,45.76,5868,0,El Cajon,1,0,Cable,32.79697,-116.969082,1,96.1,2,1,None,55277,0,0,1,0,62,1,722.0,2837.12,0.0,6019.35,0,0,92020
3625,0,0,1,0,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.85,1379.6,0,44,0,18.41,4121,0,El Cajon,0,0,NA,32.832706,-116.873258,1,19.85,0,10,None,61872,0,0,1,0,71,0,0.0,1307.11,0.0,1379.6,0,0,92021
3626,1,0,0,1,23,1,0,DSL,0,1,0,0,Month-to-month,1,Bank transfer (automatic),55.3,1284.2,0,25,47,1.58,4028,0,Encinitas,0,1,Cable,33.054579,-117.25665,0,55.3,3,0,Offer D,47126,1,0,0,1,23,0,604.0,36.34,0.0,1284.2,1,0,92024
3627,0,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,296.15,0,35,0,20.65,5052,0,Escondido,0,0,NA,33.081478000000004,-117.03381399999999,0,20.1,0,0,Offer D,49281,0,0,0,0,16,0,0.0,330.4,0.0,296.15,0,0,92025
3628,1,0,0,0,9,1,0,DSL,1,0,1,0,Month-to-month,1,Mailed check,69.5,653.25,0,24,51,34.43,3628,0,Escondido,1,1,DSL,33.21846,-117.11691599999999,0,69.5,0,0,None,43436,1,1,0,1,9,2,0.0,309.87,0.0,653.25,1,1,92026
3629,1,0,1,1,17,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,25.15,412.6,0,33,0,45.24,3931,0,Escondido,0,1,NA,33.141265000000004,-116.967221,1,25.15,3,8,Offer D,48690,0,0,1,0,17,0,0.0,769.08,0.0,412.6,0,0,92027
3630,0,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.95,85.5,1,36,0,2.01,5822,1,Fallbrook,0,0,NA,33.362575,-117.299644,0,20.95,0,0,None,42239,0,0,0,0,4,8,0.0,8.04,0.0,85.5,0,0,92028
3631,0,1,1,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.55,49.55,1,73,10,24.24,4989,1,Escondido,0,0,Fiber Optic,33.079834000000005,-117.134275,1,51.532,0,1,Offer E,17944,0,0,1,0,1,5,0.0,24.24,0.0,49.55,0,0,92029
3632,0,0,1,0,24,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,79.65,1928.7,0,24,82,44.93,3816,0,Julian,1,0,Fiber Optic,32.980678000000005,-116.262854,1,79.65,0,2,None,3577,0,0,1,1,24,1,0.0,1078.32,0.0,1928.7,1,1,92036
3633,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.25,71.25,0,68,2,17.6,5033,0,La Jolla,0,0,Fiber Optic,32.853743,-117.25034,0,71.25,0,0,None,42617,0,0,0,0,1,0,0.0,17.6,0.0,71.25,0,1,92037
3634,1,1,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),113.8,7845.8,0,75,26,24.67,4598,0,Lakeside,1,1,DSL,32.909873,-116.906774,0,113.8,0,0,None,42277,1,0,0,0,72,0,0.0,1776.2400000000002,0.0,7845.8,0,1,92040
3635,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,24.55,1750.7,0,41,0,8.98,4169,0,Oceanside,0,0,NA,33.351059,-117.420557,1,24.55,0,8,None,98239,0,0,1,0,72,2,0.0,646.5600000000002,0.0,1750.7,0,0,92054
3636,0,0,0,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.7,216.2,0,57,0,44.88,3838,0,Oceanside,0,0,NA,33.194742,-117.29032,0,19.7,1,0,Offer D,52895,0,0,0,0,11,1,0.0,493.68,0.0,216.2,0,0,92056
3637,1,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,178.5,1,37,0,8.91,3361,1,Oceanside,0,1,NA,33.254497,-117.28587900000001,0,20.25,0,0,None,46893,0,0,0,0,9,2,0.0,80.19,0.0,178.5,0,0,92057
3638,0,1,1,0,2,1,0,DSL,0,1,0,0,Month-to-month,0,Credit card (automatic),50.15,115.1,1,75,22,6.86,5461,1,Pala,0,0,Fiber Optic,33.384345,-117.07261899999999,1,52.156000000000006,0,1,Offer E,1831,0,1,1,0,2,4,25.0,13.72,0.0,115.1,0,0,92059
3639,0,1,1,0,60,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),100.5,6029,0,74,26,27.68,6442,0,Palomar Mountain,1,0,Fiber Optic,33.309852,-116.82309099999999,1,100.5,0,3,None,234,0,0,1,0,60,2,0.0,1660.8,0.0,6029.0,0,1,92060
3640,1,1,1,0,29,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,95.9,2745.2,1,70,23,35.38,2151,1,Pauma Valley,1,1,Fiber Optic,33.313828,-116.940501,1,99.736,0,1,Offer C,2615,0,0,1,1,29,6,631.0,1026.02,0.0,2745.2,0,0,92061
3641,0,0,0,0,49,1,0,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),74.45,3721.9,0,58,13,7.51,4517,0,Poway,1,0,Fiber Optic,32.984395,-117.01345400000001,0,74.45,0,0,Offer B,47969,1,0,0,1,49,1,48.38,367.99,0.0,3721.9,0,1,92064
3642,0,1,0,0,30,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.1,3121.1,0,80,21,41.93,5655,0,Ramona,1,0,Fiber Optic,33.044540999999995,-116.833922,0,104.1,0,0,None,33104,0,0,0,0,30,1,0.0,1257.9,0.0,3121.1,0,1,92065
3643,0,0,1,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.05,990.45,0,50,0,46.24,6160,0,Ranchita,0,0,NA,33.215251,-116.53633,1,19.05,0,5,Offer B,339,0,0,1,0,53,0,0.0,2450.7200000000007,0.0,990.45,0,0,92066
3644,1,0,0,1,39,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.0,1004.35,0,52,0,49.95,4295,0,Rancho Santa Fe,0,1,NA,33.012751,-117.200617,0,25.0,3,0,None,7615,0,0,0,0,39,0,0.0,1948.05,0.0,1004.35,0,0,92067
3645,0,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.05,157.65,0,45,0,31.28,3248,0,San Marcos,0,0,NA,33.162624,-117.17086299999998,0,19.05,0,0,Offer E,52664,0,0,0,0,9,0,0.0,281.52,0.0,157.65,0,0,92069
3646,1,0,0,0,39,1,0,Fiber optic,0,0,0,0,One year,0,Electronic check,81.9,3219.75,0,47,29,35.13,3446,0,Santa Ysabel,1,1,Fiber Optic,33.174725,-116.743329,0,81.9,0,0,None,1143,1,0,0,0,39,0,934.0,1370.0700000000004,0.0,3219.75,0,0,92070
3647,1,1,0,0,8,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.7,572.85,0,66,5,41.85,5242,0,Santee,0,1,Fiber Optic,32.847336,-116.99760500000001,0,69.7,0,0,Offer E,53510,0,1,0,0,8,1,29.0,334.8,0.0,572.85,0,0,92071
3648,0,0,1,1,51,1,1,Fiber optic,0,0,0,1,One year,1,Electronic check,90.15,4554.85,0,21,59,19.9,5692,0,Solana Beach,1,0,Fiber Optic,33.001813,-117.263628,1,90.15,3,4,Offer B,12173,0,2,1,1,51,2,0.0,1014.9,0.0,4554.85,1,1,92075
3649,1,0,1,1,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.35,1847.55,0,21,0,9.2,5747,0,San Marcos,0,1,NA,33.119028,-117.166036,1,25.35,2,2,None,6760,0,0,1,0,71,2,0.0,653.1999999999998,0.0,1847.55,1,0,92078
3650,1,1,0,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.65,1766.75,0,79,0,4.75,4788,0,Valley Center,0,1,NA,33.252829999999996,-116.986079,0,24.65,0,0,Offer A,14575,0,0,0,0,71,1,0.0,337.25,0.0,1766.75,0,0,92082
3651,0,1,1,0,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.55,1462.05,0,73,0,15.9,5209,0,Vista,0,0,NA,33.17494,-117.24276100000002,1,19.55,0,2,Offer A,62036,0,0,1,0,70,0,0.0,1113.0,0.0,1462.05,0,0,92083
3652,0,1,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,25.25,25.25,1,77,16,0.0,4628,1,Vista,0,0,Fiber Optic,33.22784,-117.200024,0,26.26,0,0,Offer E,44692,0,1,0,0,1,1,0.0,0.0,0.0,25.25,0,0,92084
3653,1,0,1,0,38,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),60.0,2193.2,0,47,25,0.0,2187,0,Warner Springs,0,1,Fiber Optic,33.323705,-116.626907,1,60.0,0,5,None,1205,1,0,1,1,38,0,0.0,0.0,0.0,2193.2,0,1,92086
3654,0,0,1,0,28,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Credit card (automatic),89.9,2433.5,0,56,19,33.09,3676,0,Rancho Santa Fe,1,0,Fiber Optic,32.993559999999995,-117.207121,1,89.9,0,7,None,1072,0,0,1,1,28,2,0.0,926.52,0.0,2433.5,0,1,92091
3655,0,0,1,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.4,641.15,0,57,0,12.35,3846,0,San Diego,0,0,NA,32.725229999999996,-117.171346,1,19.4,0,1,None,27505,0,0,1,0,32,0,0.0,395.2,0.0,641.15,0,0,92101
3656,1,1,1,0,49,1,0,DSL,0,1,0,0,Two year,0,Mailed check,49.8,2398.4,0,74,15,1.67,4306,0,San Diego,0,1,DSL,32.716007,-117.11746200000002,1,49.8,0,4,None,47140,0,0,1,0,49,2,35.98,81.83,0.0,2398.4,0,1,92102
3657,0,0,1,1,37,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.1,861.85,0,40,0,44.68,3753,0,San Diego,0,0,NA,32.747484,-117.166877,1,24.1,1,5,None,30202,0,0,1,0,37,0,0.0,1653.16,0.0,861.85,0,0,92103
3658,0,0,0,0,10,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,54.25,583,0,41,29,12.96,2253,0,San Diego,1,0,DSL,32.741499,-117.12740900000001,0,54.25,0,0,Offer D,47689,1,1,0,0,10,3,0.0,129.60000000000002,0.0,583.0,0,1,92104
3659,1,0,1,0,67,1,1,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),109.9,7332.4,0,36,24,23.13,5416,0,San Diego,1,1,DSL,32.741859000000005,-117.09035300000001,1,109.9,0,1,None,73006,0,0,1,1,67,0,1760.0,1549.71,0.0,7332.4,0,0,92105
3660,1,0,0,0,7,0,No phone service,DSL,0,0,0,0,One year,1,Credit card (automatic),35.5,249.55,0,28,48,0.0,5124,0,San Diego,1,1,DSL,32.71346,-117.236378,0,35.5,0,0,Offer E,18525,1,0,0,0,7,1,0.0,0.0,0.0,249.55,1,1,92106
3661,0,0,0,0,51,1,0,Fiber optic,0,0,1,1,One year,0,Credit card (automatic),87.55,4475.9,0,36,7,14.37,6021,0,San Diego,0,0,Fiber Optic,32.741852,-117.243453,0,87.55,0,0,Offer B,27959,0,0,0,1,51,1,313.0,732.87,0.0,4475.9,0,0,92107
3662,0,0,0,0,9,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.15,416.45,1,38,2,15.62,3757,1,San Diego,0,0,Cable,32.774046000000006,-117.142454,0,46.956,0,0,None,11650,0,1,0,0,9,4,0.0,140.57999999999998,0.0,416.45,0,1,92108
3663,0,0,0,0,9,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,88.4,788.6,0,23,52,35.45,2952,0,San Diego,0,0,DSL,32.787836,-117.232376,0,88.4,0,0,Offer E,46086,0,0,0,1,9,2,410.0,319.05,0.0,788.6,1,0,92109
3664,1,0,0,0,4,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.8,202.3,0,58,21,1.88,4521,0,San Diego,0,1,Cable,32.76501,-117.19938,0,50.8,0,0,Offer E,24169,1,0,0,0,4,1,0.0,7.52,0.0,202.3,0,1,92110
3665,1,0,1,0,71,1,1,Fiber optic,1,1,1,0,Two year,1,Electronic check,99.0,6994.6,0,50,6,44.06,5295,0,San Diego,1,1,Fiber Optic,32.805518,-117.16905200000001,1,99.0,0,5,None,46828,0,0,1,0,71,1,0.0,3128.26,0.0,6994.6,0,1,92111
3666,0,0,1,1,50,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),84.4,4116.15,1,59,19,35.33,5135,1,San Diego,0,0,Cable,32.697098,-117.11658700000001,1,87.77600000000002,0,1,None,47431,0,1,1,0,50,1,0.0,1766.5,0.0,4116.15,0,1,92113
3667,0,1,1,1,24,1,0,Fiber optic,0,0,1,1,Two year,1,Electronic check,96.55,2263.45,0,69,23,20.78,4309,0,San Diego,1,0,Fiber Optic,32.707892,-117.05512,1,96.55,1,9,None,66838,0,0,1,1,24,0,0.0,498.72,0.0,2263.45,0,1,92114
3668,1,0,1,0,22,1,0,DSL,1,0,1,0,One year,1,Bank transfer (automatic),59.75,1374.35,0,22,51,6.03,3947,0,San Diego,0,1,DSL,32.762506,-117.07245,1,59.75,0,10,Offer D,56887,0,0,1,0,22,0,70.09,132.66,0.0,1374.35,1,1,92115
3669,1,0,0,0,44,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,111.5,4915.15,0,48,19,44.45,2827,0,San Diego,1,1,DSL,32.765299,-117.122565,0,111.5,0,0,Offer B,33083,0,0,0,1,44,1,934.0,1955.8,0.0,4915.15,0,0,92116
3670,0,0,1,1,33,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),24.25,838.5,0,49,0,9.97,5531,0,San Diego,0,0,NA,32.825086,-117.199424,1,24.25,2,2,None,51213,0,0,1,0,33,1,0.0,329.0100000000001,0.0,838.5,0,0,92117
3671,0,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.1,75.1,1,36,9,5.94,4335,1,Coronado,0,0,Cable,32.68674,-117.18661200000001,0,78.104,0,0,None,24093,0,0,0,0,1,4,0.0,5.94,0.0,75.1,0,0,92118
3672,0,0,1,0,54,1,1,DSL,0,0,1,1,One year,1,Credit card (automatic),70.15,3715.65,1,50,13,42.1,4596,1,San Diego,0,0,DSL,32.802959,-117.02709499999999,1,72.956,0,1,None,21866,0,3,1,1,54,3,0.0,2273.4,0.0,3715.65,0,1,92119
3673,1,0,0,0,42,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.75,4273.45,1,64,18,18.79,5545,1,San Diego,0,1,DSL,32.807867,-117.060993,0,105.82,0,0,None,25569,0,0,0,1,42,0,0.0,789.18,0.0,4273.45,0,1,92120
3674,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.8,45.8,1,41,20,22.11,5973,1,San Diego,0,0,DSL,32.898613,-117.202937,0,47.632,0,0,Offer E,4258,0,1,0,0,1,5,0.0,22.11,0.0,45.8,0,0,92121
3675,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.5,20.5,0,54,0,8.56,4454,0,San Diego,0,0,NA,32.85723,-117.209774,0,20.5,0,0,None,34902,0,0,0,0,1,0,0.0,8.56,0.0,20.5,0,0,92122
3676,1,0,0,0,30,1,0,DSL,1,1,1,0,One year,0,Electronic check,70.4,2044.75,0,47,22,32.41,3380,0,San Diego,0,1,DSL,32.808814,-117.134694,0,70.4,0,0,None,25232,1,0,0,0,30,1,450.0,972.3,0.0,2044.75,0,0,92123
3677,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,30.55,30.55,0,60,9,0.0,5565,0,San Diego,0,0,Fiber Optic,32.827238,-117.08928700000001,0,30.55,0,0,None,30206,1,0,0,0,1,1,0.0,0.0,0.0,30.55,0,1,92124
3678,1,0,1,1,16,1,1,DSL,1,1,1,1,Month-to-month,0,Electronic check,84.9,1398.25,0,22,59,9.16,2269,0,San Diego,0,1,Fiber Optic,32.886925,-117.152162,1,84.9,2,5,Offer D,74232,1,0,1,1,16,0,825.0,146.56,0.0,1398.25,1,0,92126
3679,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.1,20.1,1,63,0,40.83,4933,1,San Diego,0,1,NA,33.017518,-117.11845600000001,0,20.1,0,0,Offer E,20046,0,0,0,0,1,1,0.0,40.83,0.0,20.1,0,0,92127
3680,1,0,1,0,9,0,No phone service,DSL,0,0,1,0,Month-to-month,0,Mailed check,40.65,328.95,1,64,29,0.0,4800,1,San Diego,0,1,Fiber Optic,33.000269,-117.072093,1,42.276,0,2,Offer E,42733,1,3,1,0,9,1,95.0,0.0,0.0,328.95,0,0,92128
3681,1,1,1,0,46,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.0,4680.05,1,80,24,5.36,2436,1,San Diego,1,1,Cable,32.961064,-117.13491699999999,1,105.04,0,1,Offer B,47224,0,1,1,0,46,4,1123.0,246.56,0.0,4680.05,0,0,92129
3682,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.1,69.1,1,62,20,38.66,5795,1,San Diego,0,1,Cable,32.957195,-117.202542,0,71.86399999999998,0,0,Offer E,28201,0,0,0,0,1,3,0.0,38.66,0.0,69.1,0,0,92130
3683,1,0,1,0,71,1,0,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),54.5,3778.2,0,21,59,48.32,4957,0,San Diego,0,1,Fiber Optic,32.89325,-117.08709099999999,1,54.5,0,5,None,29283,1,0,1,0,71,0,222.91,3430.72,0.0,3778.2,1,1,92131
3684,1,0,0,0,43,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.35,3161.4,0,39,28,19.66,4898,0,San Diego,0,1,DSL,32.677716,-117.04766599999999,0,75.35,0,0,Offer B,36351,0,0,0,0,43,3,0.0,845.38,0.0,3161.4,0,1,92139
3685,1,0,1,0,50,0,No phone service,DSL,1,0,1,0,One year,1,Bank transfer (automatic),44.45,2188.45,0,20,73,0.0,5363,0,San Diego,0,1,Fiber Optic,32.578103000000006,-117.012975,1,44.45,0,3,Offer B,68776,1,0,1,0,50,0,0.0,0.0,0.0,2188.45,1,1,92154
3686,0,0,0,0,13,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,75.0,999.45,1,25,53,6.03,2189,1,San Ysidro,0,0,DSL,32.555828000000005,-117.04007299999999,0,78.0,0,0,Offer D,28488,0,0,0,1,13,4,530.0,78.39,0.0,999.45,1,0,92173
3687,1,0,1,1,19,1,0,Fiber optic,0,1,1,1,One year,0,Bank transfer (automatic),100.0,1888.65,1,56,22,43.95,2608,1,Indio,0,1,Cable,33.713891,-116.237257,1,104.0,0,1,None,56307,1,0,1,1,19,0,416.0,835.0500000000002,0.0,1888.65,0,0,92201
3688,0,0,0,0,41,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),98.05,3990.6,0,43,4,29.19,5614,0,Indio,1,0,Fiber Optic,33.752938,-116.23005500000001,0,98.05,0,0,Offer B,2743,0,0,0,1,41,2,0.0,1196.79,0.0,3990.6,0,1,92203
3689,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.15,71.15,1,78,24,24.75,5287,1,Indian Wells,0,0,Fiber Optic,33.537646,-116.29108899999999,0,73.99600000000002,0,0,Offer E,3873,0,0,0,0,1,2,0.0,24.75,0.0,71.15,0,0,92210
3690,0,0,0,0,24,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Credit card (automatic),54.15,1240.25,1,25,57,0.0,5153,1,Palm Desert,1,0,Fiber Optic,33.762759,-116.324817,0,56.316,0,0,Offer C,19702,0,1,0,1,24,1,0.0,0.0,0.0,1240.25,1,1,92211
3691,0,0,1,0,40,1,1,DSL,0,1,1,0,One year,0,Bank transfer (automatic),63.9,2635,0,27,52,42.1,2654,0,Banning,0,0,Fiber Optic,33.936298,-116.849577,1,63.9,0,4,Offer B,25859,0,1,1,0,40,1,1370.0,1684.0,0.0,2635.0,1,0,92220
3692,0,0,1,1,3,1,1,DSL,0,1,1,0,Month-to-month,1,Bank transfer (automatic),69.15,235,0,23,73,24.28,2301,0,Beaumont,1,0,Fiber Optic,33.946982,-116.977672,1,69.15,3,3,None,17721,0,0,1,0,3,4,172.0,72.84,0.0,235.0,1,0,92223
3693,0,0,0,0,37,1,1,DSL,1,0,1,0,One year,0,Bank transfer (automatic),64.65,2347.85,0,42,9,37.18,5255,0,Blythe,0,0,Fiber Optic,33.674583,-114.71611999999999,0,64.65,0,0,None,24659,0,0,0,0,37,0,211.0,1375.66,0.0,2347.85,0,0,92225
3694,0,0,1,1,67,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),108.75,7156.2,1,59,31,32.15,5516,1,Brawley,1,0,Cable,33.03933,-115.19185700000001,1,113.1,0,1,None,23394,1,3,1,1,67,1,2218.0,2154.05,0.0,7156.2,0,0,92227
3695,0,0,1,1,32,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,98.85,3089.6,0,59,22,24.04,3149,0,Cabazon,0,0,DSL,33.929812,-116.76058,1,98.85,1,2,None,2355,0,0,1,1,32,0,0.0,769.28,0.0,3089.6,0,1,92230
3696,0,0,1,0,6,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.15,270.8,1,59,31,6.94,5271,1,Calexico,0,0,Cable,32.690653999999995,-115.431225,1,51.11600000000001,0,1,Offer E,27804,1,0,1,0,6,0,84.0,41.64,0.0,270.8,0,0,92231
3697,0,0,1,1,32,1,1,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,89.6,2901.8,0,25,82,48.49,4444,0,Calipatria,0,0,Fiber Optic,33.143826000000004,-115.49748500000001,1,89.6,3,6,None,7857,0,2,1,0,32,1,2379.0,1551.68,0.0,2901.8,1,0,92233
3698,0,0,0,0,59,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,83.25,4949.1,0,48,16,31.23,4094,0,Cathedral City,1,0,Fiber Optic,33.829583,-116.474131,0,83.25,0,0,Offer B,43141,0,0,0,0,59,0,792.0,1842.57,0.0,4949.1,0,0,92234
3699,0,0,1,0,30,1,0,DSL,0,1,0,1,One year,0,Bank transfer (automatic),70.25,2198.9,0,53,13,17.33,5417,0,Coachella,1,0,Fiber Optic,33.680031,-116.171678,1,70.25,0,7,None,23170,1,0,1,1,30,0,0.0,519.9,0.0,2198.9,0,1,92236
3700,1,0,0,1,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.4,374.5,1,30,0,22.78,3785,1,Desert Center,0,1,NA,33.889604999999996,-115.25700900000001,0,19.4,3,0,None,964,0,0,0,0,20,4,0.0,455.6,0.0,374.5,0,0,92239
3701,0,0,1,1,27,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,24.5,761.95,0,51,0,35.52,2645,0,Desert Hot Springs,0,0,NA,33.948558,-116.516976,1,24.5,1,1,None,22796,0,1,1,0,27,3,0.0,959.04,0.0,761.95,0,0,92240
3702,0,1,0,0,20,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,79.15,1520.9,1,69,6,11.82,4997,1,Desert Hot Springs,0,0,Fiber Optic,33.832799,-116.250973,0,82.316,0,0,None,5529,0,0,0,0,20,4,91.0,236.4,0.0,1520.9,0,0,92241
3703,1,0,0,1,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,190.25,0,60,0,27.34,3444,0,Earp,0,1,NA,34.137741999999996,-114.36514,0,20.1,3,0,None,1564,0,0,0,0,9,2,0.0,246.06,0.0,190.25,0,0,92242
3704,0,0,1,1,68,1,1,DSL,1,1,1,0,One year,1,Credit card (automatic),73.0,5163,0,47,16,20.15,4156,0,El Centro,1,0,Fiber Optic,32.770393,-115.60915,1,73.0,2,8,None,43712,0,0,1,0,68,2,826.0,1370.1999999999996,0.0,5163.0,0,0,92243
3705,0,0,1,1,69,1,1,DSL,1,0,0,0,Two year,0,Credit card (automatic),61.4,4059.85,0,56,19,39.07,5266,0,Heber,0,0,Fiber Optic,32.730583,-115.50108300000001,1,61.4,2,10,None,3535,1,0,1,0,69,1,771.0,2695.83,0.0,4059.85,0,0,92249
3706,1,0,0,0,26,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,84.3,2281.6,0,62,30,37.69,5471,0,Holtville,1,1,Fiber Optic,32.811001,-115.15286499999999,0,84.3,0,0,None,8062,1,0,0,0,26,1,684.0,979.94,0.0,2281.6,0,0,92250
3707,1,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.9,1356.7,0,49,0,28.19,6058,0,Imperial,0,1,NA,32.858595,-115.662709,1,19.9,2,10,Offer A,14546,0,0,1,0,69,1,0.0,1945.11,0.0,1356.7,0,0,92251
3708,1,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.4,231.45,0,60,0,49.8,5397,0,Joshua Tree,0,1,NA,34.167235999999995,-116.28151100000001,0,20.4,0,0,Offer D,8141,0,0,0,0,11,1,0.0,547.8,0.0,231.45,0,0,92252
3709,1,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.75,50.75,0,19,26,24.66,3631,0,La Quinta,0,1,DSL,33.695532,-116.310571,0,50.75,0,0,None,23971,0,0,0,0,1,1,0.0,24.66,0.0,50.75,1,1,92253
3710,1,0,1,1,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.45,242.4,0,37,0,37.59,4613,0,Mecca,0,1,NA,33.543834999999994,-115.99390600000001,1,20.45,1,0,Offer D,8768,0,0,0,0,10,2,0.0,375.9,0.0,242.4,0,0,92254
3711,0,0,1,1,55,1,1,DSL,1,1,0,1,One year,1,Bank transfer (automatic),75.75,4264.25,0,41,29,16.16,4489,0,Morongo Valley,0,0,DSL,34.097863000000004,-116.59456100000001,1,75.75,3,7,Offer B,3499,1,0,1,1,55,0,0.0,888.8,0.0,4264.25,0,1,92256
3712,1,0,0,0,44,1,0,DSL,1,0,1,0,One year,0,Electronic check,65.4,2774.55,0,42,2,34.98,5827,0,Niland,0,1,Fiber Optic,33.345825,-115.596574,0,65.4,0,0,Offer B,2753,1,0,0,0,44,0,55.0,1539.12,0.0,2774.55,0,0,92257
3713,1,1,1,0,46,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.4,3605.2,1,71,3,48.62,4876,1,North Palm Springs,0,1,DSL,33.906496000000004,-116.569499,1,83.61600000000001,0,1,Offer B,732,0,0,1,0,46,2,108.0,2236.52,0.0,3605.2,0,0,92258
3714,1,0,1,1,69,1,0,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),59.75,4069.9,0,32,12,49.4,4665,0,Ocotillo,1,1,DSL,32.698964000000004,-115.886656,1,59.75,1,4,Offer A,471,0,0,1,0,69,0,0.0,3408.6,0.0,4069.9,0,1,92259
3715,1,1,0,0,11,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,78.5,874.2,0,71,3,41.58,4333,0,Palm Desert,0,1,Fiber Optic,33.694501,-116.41271100000002,0,78.5,0,0,None,29340,0,0,0,1,11,1,26.0,457.38,0.0,874.2,0,0,92260
3716,0,0,1,0,11,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,102.0,1145.35,1,36,11,7.89,5750,1,Palm Springs,0,0,Fiber Optic,33.839989,-116.65921499999999,1,106.08,0,1,None,24924,0,1,1,1,11,2,0.0,86.78999999999998,0.0,1145.35,0,1,92262
3717,1,0,0,0,29,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),48.95,1323.7,0,34,25,10.06,4825,0,Palm Springs,1,1,Fiber Optic,33.745746000000004,-116.514215,0,48.95,0,0,Offer C,18884,0,0,0,0,29,0,33.09,291.74,0.0,1323.7,0,1,92264
3718,0,0,1,0,57,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,99.65,5497.05,0,32,16,12.19,5106,0,Palo Verde,0,0,Cable,33.3249,-114.758334,1,99.65,0,0,Offer B,291,0,1,0,1,57,2,0.0,694.8299999999998,0.0,5497.05,0,1,92266
3719,1,0,0,0,28,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),18.25,534.7,0,58,0,40.39,5327,0,Parker Dam,0,1,NA,34.273872,-114.192901,0,18.25,0,0,Offer C,131,0,0,0,0,28,0,0.0,1130.92,0.0,534.7,0,0,92267
3720,0,0,0,0,42,1,0,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),54.55,2455.05,0,42,8,32.16,5387,0,Pioneertown,1,0,Cable,34.201108000000005,-116.593456,0,54.55,0,0,Offer B,354,0,0,0,0,42,1,0.0,1350.7199999999998,0.0,2455.05,0,1,92268
3721,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.65,38.7,1,60,0,24.71,3845,1,Rancho Mirage,0,0,NA,33.763678000000006,-116.429928,0,20.65,0,0,Offer E,12465,0,0,0,0,2,5,0.0,49.42,0.0,38.7,0,0,92270
3722,1,0,0,1,23,0,No phone service,DSL,1,1,0,0,One year,0,Bank transfer (automatic),40.65,947.4,0,61,19,0.0,5230,0,Seeley,0,1,Cable,32.790282,-115.689559,0,40.65,1,0,None,1632,1,0,0,0,23,1,180.0,0.0,0.0,947.4,0,0,92273
3723,0,0,1,1,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.45,357,0,39,0,14.6,2047,0,Thermal,0,0,NA,33.53604,-116.119222,1,20.45,2,8,None,17018,0,0,1,0,18,0,0.0,262.8,0.0,357.0,0,0,92274
3724,1,0,1,1,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),24.8,1476.25,0,60,0,16.48,5105,0,Salton City,0,1,NA,33.28156,-115.955541,1,24.8,1,1,None,799,0,0,1,0,62,0,0.0,1021.76,0.0,1476.25,0,0,92275
3725,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.8,70.8,1,23,30,30.6,3901,1,Thousand Palms,0,0,Cable,33.849263,-116.382778,0,73.632,0,0,Offer E,6242,0,0,0,1,1,2,0.0,30.6,0.0,70.8,1,0,92276
3726,1,0,0,0,16,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),89.05,1448.6,1,37,20,11.96,5953,1,Escondido,0,1,Cable,33.141265000000004,-116.967221,0,92.61200000000001,0,0,None,48690,1,0,0,1,16,0,290.0,191.36,0.0,1448.6,0,0,92027
3727,0,0,0,0,3,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.6,291.9,1,48,14,9.95,3260,1,Twentynine Palms,0,0,Cable,34.457829,-116.13958899999999,0,100.464,0,0,Offer E,14104,0,1,0,1,3,3,4.09,29.85,0.0,291.9,0,1,92278
3728,1,0,0,0,67,1,1,DSL,1,1,1,1,One year,1,Bank transfer (automatic),88.8,5903.15,0,19,59,37.32,4081,0,Escondido,1,1,DSL,33.141265000000004,-116.967221,0,88.8,0,0,Offer A,48690,1,0,0,1,67,0,3483.0,2500.44,0.0,5903.15,1,0,92027
3729,1,0,0,0,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.05,1201.65,0,19,0,33.68,4568,0,Westmorland,0,1,NA,33.03679,-115.60503,0,20.05,0,0,None,2388,0,0,0,0,62,1,0.0,2088.16,0.0,1201.65,1,0,92281
3730,0,0,1,0,57,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),104.5,5921.35,1,47,28,40.13,4471,1,White Water,1,0,Cable,33.972293,-116.654195,1,108.68,0,1,None,805,0,2,1,1,57,1,1658.0,2287.4100000000008,0.0,5921.35,0,0,92282
3731,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.8,146.65,0,31,14,11.19,3527,0,Winterhaven,0,1,DSL,32.852947,-114.850784,0,69.8,0,0,None,3663,0,0,0,0,2,0,21.0,22.38,0.0,146.65,0,0,92283
3732,0,0,1,1,23,1,1,DSL,1,0,1,0,Two year,1,Bank transfer (automatic),77.15,1759.4,0,62,12,33.02,2572,0,Yucca Valley,1,0,Fiber Optic,34.159534,-116.42598400000001,1,77.15,2,10,None,20486,1,0,1,0,23,1,0.0,759.46,0.0,1759.4,0,1,92284
3733,0,0,0,1,25,0,No phone service,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),35.05,844.45,0,32,75,0.0,2754,0,Landers,0,0,DSL,34.341737,-116.53941599999999,0,35.05,3,0,Offer C,2182,1,0,0,0,25,0,0.0,0.0,0.0,844.45,0,1,92285
3734,0,1,0,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),108.1,7774.05,0,65,20,26.87,4474,0,Adelanto,1,0,Fiber Optic,34.667815000000004,-117.53618300000001,0,108.1,0,0,Offer A,18980,1,0,0,1,72,1,0.0,1934.64,0.0,7774.05,0,1,92301
3735,0,0,1,0,2,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.05,134.05,0,40,13,22.23,2115,0,Amboy,0,0,Fiber Optic,34.559882,-115.63716399999998,1,84.05,0,9,None,42,0,0,1,0,2,2,0.0,44.46,0.0,134.05,0,1,92304
3736,0,0,0,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.2,140.95,0,26,0,5.27,5066,0,Angelus Oaks,0,0,NA,34.1678,-116.86433000000001,0,20.2,0,0,None,301,0,0,0,0,8,0,0.0,42.16,0.0,140.95,1,0,92305
3737,0,0,0,0,5,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.6,249.95,1,54,2,37.1,2353,1,Fallbrook,0,0,DSL,33.362575,-117.299644,0,52.623999999999995,0,0,Offer E,42239,0,0,0,0,5,0,5.0,185.5,0.0,249.95,0,0,92028
3738,1,0,0,0,35,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Electronic check,49.2,1701.65,0,47,26,0.0,2782,0,Apple Valley,1,1,DSL,34.424926,-117.184503,0,49.2,0,0,Offer C,28819,0,0,0,1,35,0,0.0,0.0,0.0,1701.65,0,1,92308
3739,1,0,0,0,24,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,24.6,592.65,0,60,0,47.33,5448,0,Baker,0,1,NA,35.28952,-116.09221399999998,0,24.6,0,0,Offer C,904,0,0,0,0,24,2,0.0,1135.92,0.0,592.65,0,0,92309
3740,0,0,1,1,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.65,135.75,0,33,10,29.03,3916,0,Fort Irwin,0,0,Cable,35.349241,-116.77028100000001,1,71.65,1,5,None,9465,0,0,1,0,2,0,0.0,58.06,0.0,135.75,0,1,92310
3741,1,0,1,1,72,1,1,Fiber optic,1,1,0,1,Two year,1,Credit card (automatic),104.9,7732.65,0,38,25,32.22,6378,0,Barstow,1,1,DSL,34.965648,-117.00150900000001,1,104.9,3,6,Offer A,31293,1,0,1,1,72,0,0.0,2319.84,0.0,7732.65,0,1,92311
3742,0,0,0,0,41,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,106.5,4282.4,0,20,59,36.7,4434,0,Grand Terrace,1,0,Fiber Optic,34.029175,-117.30721100000001,0,106.5,0,0,None,11024,1,0,0,0,41,0,0.0,1504.7,0.0,4282.4,1,1,92313
3743,1,0,0,1,4,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,49.35,219.65,1,40,30,26.04,5858,1,Big Bear City,0,1,Cable,34.278967,-116.773825,0,51.32400000000001,1,0,Offer E,9899,0,1,0,0,4,4,0.0,104.16,0.0,219.65,0,1,92314
3744,1,0,0,0,26,1,0,Fiber optic,0,1,0,0,One year,0,Bank transfer (automatic),75.5,2018.1,0,59,29,39.63,5184,0,Big Bear Lake,0,1,Fiber Optic,34.242058,-116.89801999999999,0,75.5,0,0,Offer C,5447,0,0,0,0,26,0,585.0,1030.38,0.0,2018.1,0,0,92315
3745,1,0,0,0,7,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,94.25,669,1,22,76,12.05,5267,1,Bloomington,0,1,DSL,34.059722,-117.39103999999999,0,98.02,0,0,Offer E,25995,0,4,0,1,7,5,508.0,84.35000000000002,0.0,669.0,1,0,92316
3746,0,0,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,68.95,68.95,1,64,14,21.65,5644,1,Calimesa,0,0,DSL,33.982787,-117.057627,1,71.708,0,1,Offer E,7334,0,1,1,0,1,3,0.0,21.65,0.0,68.95,0,0,92320
3747,0,0,1,1,4,1,1,DSL,0,1,0,0,Month-to-month,1,Mailed check,58.5,224.85,0,28,52,35.2,5605,0,Cedar Glen,0,0,Cable,34.255203,-117.17565400000001,1,58.5,3,9,None,455,1,2,1,0,4,2,0.0,140.8,0.0,224.85,1,1,92321
3748,1,0,0,0,48,1,0,DSL,0,1,1,1,Two year,0,Credit card (automatic),78.9,3771.5,0,45,10,3.59,4063,0,Colton,1,1,Fiber Optic,34.030915,-117.273201,0,78.9,0,0,None,52202,1,0,0,1,48,2,377.0,172.32,0.0,3771.5,0,0,92324
3749,1,1,0,0,2,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.85,196.75,1,70,15,25.19,4998,1,Crestline,0,1,Cable,34.248061,-117.29028000000001,0,97.604,0,0,None,10484,0,2,0,0,2,3,30.0,50.38,0.0,196.75,0,0,92325
3750,0,1,1,0,12,1,0,DSL,1,0,1,1,One year,1,Electronic check,79.2,943.85,0,73,13,37.15,3355,0,Daggett,1,0,Fiber Optic,34.875144,-116.821698,1,79.2,0,3,None,678,1,0,1,1,12,0,0.0,445.8,0.0,943.85,0,1,92327
3751,1,0,1,0,60,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),109.45,6572.85,0,36,9,4.59,4350,0,Death Valley,1,1,Cable,36.27688,-117.033326,1,109.45,0,6,None,443,1,0,1,1,60,0,0.0,275.4,0.0,6572.85,0,1,92328
3752,1,0,0,0,55,1,0,DSL,1,0,0,0,Two year,1,Electronic check,59.2,3175.85,0,20,48,12.28,5162,0,Essex,1,1,Fiber Optic,34.9436,-115.287901,0,59.2,0,0,None,115,1,0,0,0,55,0,152.44,675.4,0.0,3175.85,1,1,92332
3753,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,29.15,29.15,0,34,22,0.0,3923,0,Fawnskin,0,1,DSL,34.274846000000004,-116.93758100000001,0,29.15,0,0,None,414,1,0,0,0,1,0,0.0,0.0,0.0,29.15,0,0,92333
3754,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,20.05,0,30,0,11.1,2313,0,Fontana,0,1,NA,34.087558,-117.464096,0,20.05,0,0,None,82630,0,0,0,0,1,1,0.0,11.1,0.0,20.05,0,0,92335
3755,1,0,0,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.05,318.9,1,62,32,42.44,3685,1,Fontana,0,1,DSL,34.136367,-117.460803,0,79.092,0,0,None,54586,0,2,0,0,4,2,0.0,169.76,0.0,318.9,0,1,92336
3756,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,24.45,24.45,1,44,2,0.0,2121,1,Fontana,0,1,Fiber Optic,34.049671000000004,-117.468896,0,25.428,0,0,None,29847,0,0,0,0,1,0,0.0,0.0,0.0,24.45,0,1,92337
3757,0,0,0,0,42,1,0,DSL,0,0,0,1,Two year,0,Credit card (automatic),66.5,2762.75,0,33,20,34.76,4668,0,Ludlow,1,0,Fiber Optic,34.702766,-116.093376,0,66.5,0,0,None,23,1,0,0,1,42,0,0.0,1459.9199999999996,0.0,2762.75,0,1,92338
3758,0,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),49.55,49.55,0,45,15,10.83,5277,0,Forest Falls,0,0,Fiber Optic,34.067699,-116.90389099999999,0,49.55,0,0,None,958,0,0,0,0,1,0,0.0,10.83,0.0,49.55,0,1,92339
3759,1,0,0,0,7,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),89.35,631.85,1,35,19,36.84,4154,1,Green Valley Lake,1,1,Cable,34.244411,-117.072654,0,92.924,0,0,None,317,0,2,0,0,7,7,120.0,257.88,0.0,631.85,0,0,92341
3760,1,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),73.6,232.5,0,29,71,27.34,5510,0,Helendale,1,1,Fiber Optic,34.757783,-117.33997,0,73.6,0,0,None,4948,0,0,0,0,3,1,16.51,82.02,0.0,232.5,1,1,92342
3761,0,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),82.65,5919.35,0,53,11,17.28,4324,0,Hesperia,1,0,Cable,34.361387,-117.33750900000001,1,82.65,0,7,Offer A,68515,0,0,1,1,72,0,65.11,1244.16,0.0,5919.35,0,1,92345
3762,1,0,0,0,15,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.0,749.25,0,40,28,11.75,2597,0,Highland,0,1,Fiber Optic,34.129677,-117.15427700000001,0,49.0,0,0,None,48245,0,0,0,0,15,0,210.0,176.25,0.0,749.25,0,0,92346
3763,1,0,1,0,4,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.35,307.4,1,60,14,32.43,4167,1,Hinkley,0,1,Cable,34.983808,-117.239306,1,83.564,0,3,None,1933,0,3,1,0,4,3,43.0,129.72,0.0,307.4,0,0,92347
3764,0,0,0,0,11,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,25.2,245.15,0,50,0,1.87,4998,0,Lake Arrowhead,0,0,NA,34.2565,-117.19335,0,25.2,0,0,None,9793,0,0,0,0,11,0,0.0,20.57,0.0,245.15,0,0,92352
3765,0,0,0,0,5,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,25.45,134.75,0,63,0,5.41,4855,0,Loma Linda,0,0,NA,34.049315,-117.255974,0,25.45,0,0,None,18068,0,0,0,0,5,1,0.0,27.05,0.0,134.75,0,0,92354
3766,0,1,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,55.8,55.8,1,66,24,26.22,5527,1,Lucerne Valley,1,0,Cable,34.508417,-116.856103,0,58.032,0,0,Offer E,5256,0,2,0,0,1,1,0.0,26.22,0.0,55.8,0,0,92356
3767,1,0,1,0,72,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),110.9,8240.85,0,37,14,46.16,4938,0,Lytle Creek,1,1,DSL,34.238162,-117.534306,1,110.9,0,6,Offer A,1090,1,0,1,1,72,1,1154.0,3323.5199999999995,0.0,8240.85,0,0,92358
3768,0,0,1,0,55,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),77.75,4266.4,0,20,53,23.45,4621,0,Mentone,0,0,Fiber Optic,34.103578000000006,-117.04054,1,77.75,0,3,None,7324,0,0,1,0,55,2,2261.0,1289.75,0.0,4266.4,1,0,92359
3769,0,0,1,1,40,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,26.2,1077.5,0,49,0,49.22,2211,0,Needles,0,0,NA,34.711224,-114.702256,1,26.2,4,5,None,5488,0,0,1,0,40,0,0.0,1968.8,0.0,1077.5,0,0,92363
3770,0,0,1,0,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.9,1115.6,0,43,0,44.86,4408,0,Nipton,0,0,NA,35.478736,-115.51698400000001,1,19.9,0,6,None,162,0,0,1,0,57,0,0.0,2557.02,0.0,1115.6,0,0,92364
3771,1,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.05,79.05,1,24,57,31.34,3555,1,Temecula,0,1,Cable,33.507255,-117.029473,0,82.212,0,0,None,46171,0,1,0,1,1,1,0.0,31.34,0.0,79.05,1,0,92592
3772,1,0,1,0,1,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,95.0,95,1,42,6,12.04,4489,1,Oro Grande,0,1,Fiber Optic,34.647959,-117.296957,1,98.8,0,1,None,909,0,3,1,1,1,3,0.0,12.04,0.0,95.0,0,0,92368
3773,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,25.2,25.2,1,29,80,0.0,3196,1,Phelan,0,0,Cable,34.441123,-117.53788600000001,0,26.208000000000002,0,0,None,12463,0,0,0,1,1,4,0.0,0.0,0.0,25.2,1,1,92371
3774,1,1,1,1,52,1,1,DSL,0,1,1,1,One year,1,Electronic check,80.85,4079.55,0,72,22,7.04,6090,0,Pinon Hills,1,1,Cable,34.459322,-117.629729,1,80.85,1,1,None,4280,0,0,1,1,52,1,0.0,366.08,0.0,4079.55,0,1,92372
3775,1,1,0,0,41,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.4,4187.75,1,77,23,42.06,2169,1,Redlands,1,1,Cable,34.003243,-117.13828600000001,0,102.336,0,0,Offer B,31230,0,0,0,0,41,0,963.0,1724.46,0.0,4187.75,0,0,92373
3776,1,0,1,0,43,1,0,DSL,0,0,1,0,One year,1,Mailed check,56.35,2391.15,0,50,23,4.34,4928,0,Redlands,0,1,DSL,34.064073,-117.16615800000001,1,56.35,0,9,None,36675,0,0,1,0,43,1,0.0,186.62,0.0,2391.15,0,1,92374
3777,0,0,1,1,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.3,890.5,0,24,0,2.56,5829,0,Rialto,0,0,NA,34.109775,-117.378904,1,19.3,3,1,None,75882,0,0,1,0,47,0,0.0,120.32,0.0,890.5,1,0,92376
3778,1,0,0,0,3,1,1,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),50.4,137.25,0,28,59,29.74,4639,0,Rialto,0,1,Cable,34.156758,-117.40468600000001,0,50.4,0,0,None,18518,0,0,0,0,3,2,81.0,89.22,0.0,137.25,1,0,92377
3779,1,1,1,1,66,1,1,DSL,1,1,1,0,Two year,0,Credit card (automatic),79.4,5154.6,1,71,16,30.03,5910,1,Running Springs,1,1,Fiber Optic,34.186211,-117.07683,1,82.57600000000002,0,1,None,5395,1,0,1,0,66,5,825.0,1981.98,0.0,5154.6,0,0,92382
3780,1,0,1,1,55,1,0,DSL,0,0,0,0,Two year,1,Credit card (automatic),55.25,3119.9,0,24,30,46.61,5821,0,Shoshone,1,1,Fiber Optic,35.924252,-116.18866799999999,1,55.25,1,5,None,87,1,0,1,0,55,2,936.0,2563.55,0.0,3119.9,1,0,92384
3781,1,0,0,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.1,529.5,0,40,0,49.52,5880,0,Sugarloaf,0,1,NA,34.243088,-116.83001499999999,0,19.1,0,0,Offer C,1834,0,0,0,0,29,1,0.0,1436.0800000000004,0.0,529.5,0,0,92386
3782,0,0,0,1,12,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.05,966.55,0,56,19,17.85,4621,0,Fallbrook,0,0,Fiber Optic,33.362575,-117.299644,0,84.05,1,0,None,42239,0,0,0,0,12,1,184.0,214.2,0.0,966.55,0,0,92028
3783,0,0,1,0,66,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.2,6936.85,0,39,30,42.23,4016,0,Victorville,1,0,DSL,34.486835,-117.362274,1,105.2,0,6,Offer A,63235,0,0,1,1,66,0,2081.0,2787.18,0.0,6936.85,0,0,92392
3784,1,1,0,0,35,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.4,3496.3,1,68,28,39.69,3689,1,Victorville,1,1,Fiber Optic,34.567058,-117.362329,0,105.456,0,0,Offer C,12083,0,0,0,0,35,0,979.0,1389.15,0.0,3496.3,0,0,92394
3785,1,1,1,0,10,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.8,914.3,1,71,26,16.88,5124,1,Wrightwood,1,1,Cable,34.358321000000004,-117.61826299999998,1,93.39200000000001,0,0,None,4253,0,0,0,0,10,3,238.0,168.79999999999995,0.0,914.3,0,0,92397
3786,1,0,1,1,27,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.75,1929,0,60,23,25.26,4994,0,Yermo,0,1,Fiber Optic,35.013298999999996,-116.834092,1,75.75,3,7,Offer C,1195,0,0,1,0,27,1,0.0,682.0200000000002,0.0,1929.0,0,1,92398
3787,0,0,0,0,58,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.3,5817.7,0,20,73,35.55,6460,0,Yucaipa,0,0,Fiber Optic,34.045970000000004,-117.011825,0,95.3,0,0,None,41575,1,0,0,1,58,0,0.0,2061.9,0.0,5817.7,1,1,92399
3788,1,0,1,0,54,1,0,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),109.75,6110.2,1,34,10,42.09,6274,1,San Bernardino,1,1,Cable,34.105934999999995,-117.2914,1,114.14,0,1,None,1779,1,0,1,1,54,0,611.0,2272.86,0.0,6110.2,0,0,92401
3789,1,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,178.8,0,56,0,40.74,2788,0,San Bernardino,0,1,NA,34.183285999999995,-117.221722,0,19.85,0,0,None,53636,0,0,0,0,9,2,0.0,366.66,0.0,178.8,0,0,92404
3790,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.3,28.3,1,56,0,15.79,2279,1,San Bernardino,0,1,NA,34.142747,-117.30086399999999,0,19.3,0,0,None,24644,0,0,0,0,2,0,0.0,31.58,0.0,28.3,0,0,92405
3791,1,0,0,0,6,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.1,435,0,59,18,18.65,5741,0,San Bernardino,0,1,Cable,34.250069,-117.39394899999999,0,69.1,0,0,Offer E,49355,0,0,0,0,6,1,0.0,111.9,0.0,435.0,0,1,92407
3792,0,1,0,0,26,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,91.25,2351.8,1,79,30,34.69,5154,1,San Bernardino,0,0,Cable,34.084909,-117.25810700000001,0,94.9,0,0,Offer C,12149,0,2,0,0,26,7,706.0,901.94,0.0,2351.8,0,0,92408
3793,0,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,186.15,0,57,0,2.6,5546,0,San Bernardino,0,0,NA,34.106922,-117.29755300000001,0,20.25,0,0,Offer E,44556,0,0,0,0,9,0,0.0,23.4,0.0,186.15,0,0,92410
3794,1,0,1,0,8,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,54.75,445.85,0,36,8,19.0,4099,0,San Bernardino,1,1,Fiber Optic,34.122501,-117.32013799999999,1,54.75,0,10,Offer E,23146,0,0,1,0,8,0,0.0,152.0,0.0,445.85,0,1,92411
3795,1,0,0,0,12,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,81.45,912,0,32,16,11.04,2916,0,Riverside,0,1,Cable,33.994676,-117.372498,0,81.45,0,0,None,18999,0,0,0,0,12,0,146.0,132.48,0.0,912.0,0,0,92501
3796,0,0,0,0,15,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.1,679.55,1,33,29,9.71,5209,1,Riverside,0,0,Cable,33.890046000000005,-117.455583,0,51.06399999999999,0,0,None,71678,0,2,0,0,15,4,197.0,145.65,0.0,679.55,0,0,92503
3797,1,0,1,0,43,1,1,DSL,1,0,1,1,One year,1,Electronic check,80.2,3581.6,0,30,69,33.97,5888,0,Riverside,1,1,DSL,33.9108,-117.39815300000001,1,80.2,0,7,None,46550,0,0,1,1,43,1,247.13,1460.71,0.0,3581.6,0,1,92504
3798,1,0,0,0,42,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.3,4222.95,0,48,13,25.69,3286,0,Riverside,0,1,Fiber Optic,33.920907,-117.489426,0,100.3,0,0,None,38446,1,0,0,1,42,0,549.0,1078.98,0.0,4222.95,0,0,92505
3799,0,0,0,0,31,1,1,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),65.25,1994.3,1,29,57,31.14,4403,1,Riverside,1,0,Fiber Optic,33.930931,-117.36178799999999,0,67.86,0,0,Offer C,42425,1,0,0,0,31,0,1137.0,965.34,0.0,1994.3,1,0,92506
3800,0,0,0,1,66,1,1,Fiber optic,1,0,0,0,Two year,1,Credit card (automatic),90.95,5930.05,0,20,51,27.09,6204,0,Riverside,1,0,Fiber Optic,33.976328,-117.31978600000001,0,90.95,1,0,Offer A,48649,1,0,0,0,66,0,0.0,1787.94,0.0,5930.05,1,1,92507
3801,0,1,0,0,18,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,85.45,1505.85,1,80,23,2.36,5145,1,Riverside,0,0,Cable,33.885498999999996,-117.324959,0,88.86800000000002,0,0,None,17147,1,0,0,0,18,3,346.0,42.48,0.0,1505.85,0,0,92508
3802,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,20,0,55,0,25.99,5650,0,Riverside,0,1,NA,34.004379,-117.447864,0,20.0,0,0,Offer E,63999,0,0,0,0,1,3,0.0,25.99,0.0,20.0,0,0,92509
3803,1,0,1,0,61,1,1,Fiber optic,0,1,1,0,Two year,1,Electronic check,94.1,5638.3,1,46,12,26.94,6295,1,March Air Reserve Base,0,1,DSL,33.888323,-117.277533,1,97.86399999999999,0,9,Offer B,1005,1,1,1,0,61,3,677.0,1643.34,0.0,5638.3,0,0,92518
3804,1,0,0,0,10,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,79.85,797.25,0,43,22,15.6,5739,0,Lake Elsinore,0,1,DSL,33.655421000000004,-117.391751,0,79.85,0,0,None,38519,0,0,0,0,10,2,0.0,156.0,0.0,797.25,0,1,92530
3805,1,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.65,71.65,1,65,13,28.46,5674,1,Lake Elsinore,0,1,DSL,33.705836,-117.31820400000001,0,74.516,0,0,Offer E,4546,0,0,0,0,1,0,0.0,28.46,0.0,71.65,0,1,92532
3806,0,1,0,0,18,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,73.55,1359.45,0,71,24,7.51,5313,0,Aguanga,0,0,Fiber Optic,33.482243,-116.827173,0,73.55,0,0,None,2433,0,0,0,0,18,0,326.0,135.18,0.0,1359.45,0,0,92536
3807,1,0,1,0,24,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.65,2542.45,1,51,16,3.0,4734,1,Anza,1,1,Cable,33.527605,-116.666551,1,108.836,0,2,Offer C,3745,0,1,1,1,24,4,407.0,72.0,0.0,2542.45,0,0,92539
3808,0,0,1,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.3,54.7,0,53,0,10.13,5722,0,Hemet,0,0,NA,33.739415,-116.96833899999999,1,19.3,2,5,None,29687,0,0,1,0,3,1,0.0,30.39,0.0,54.7,0,0,92543
3809,1,0,0,0,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.15,989.05,0,24,0,21.72,5249,0,Hemet,0,1,NA,33.644585,-116.871544,0,20.15,0,0,None,39264,0,1,0,0,50,2,0.0,1086.0,0.0,989.05,1,0,92544
3810,1,0,1,1,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.55,44.55,0,48,18,41.1,3408,0,Hemet,0,1,Fiber Optic,33.734933000000005,-117.044145,1,44.55,2,1,None,25694,0,0,1,0,1,1,0.0,41.1,0.0,44.55,0,0,92545
3811,1,0,0,0,2,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,54.45,87.3,0,32,19,19.87,5753,0,Homeland,0,1,Fiber Optic,33.761894,-117.12086799999999,0,54.45,0,0,None,4283,1,0,0,0,2,0,0.0,39.74,0.0,87.3,0,1,92548
3812,1,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.65,351.55,0,27,0,47.79,4774,0,Idyllwild,0,1,NA,33.755039000000004,-116.741796,0,19.65,0,0,None,3588,0,0,0,0,17,0,0.0,812.43,0.0,351.55,1,0,92549
3813,1,0,1,1,69,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,105.0,7297.75,0,47,11,22.49,5436,0,Moreno Valley,1,1,Fiber Optic,33.882740000000005,-117.224878,1,105.0,2,9,Offer A,22983,0,0,1,1,69,1,803.0,1551.81,0.0,7297.75,0,0,92551
3814,1,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),88.7,6301.7,0,63,19,47.66,5764,0,Moreno Valley,1,1,Fiber Optic,33.923149,-117.244933,1,88.7,0,4,Offer A,61205,1,0,1,1,72,0,0.0,3431.5199999999995,0.0,6301.7,0,1,92553
3815,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.25,210.3,1,44,30,35.54,3207,1,Moreno Valley,0,0,Cable,33.907361,-117.109972,0,77.22,0,0,None,12743,0,0,0,0,3,1,0.0,106.62,0.0,210.3,0,1,92555
3816,1,1,1,1,50,1,1,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),75.15,3822.45,0,74,18,32.9,6084,0,Moreno Valley,1,1,Fiber Optic,33.970661,-117.255039,1,75.15,2,3,None,46214,0,0,1,1,50,0,688.0,1645.0,0.0,3822.45,0,0,92557
3817,0,0,0,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.25,1048.45,0,28,0,28.46,4218,0,Mountain Center,0,0,NA,33.638645000000004,-116.55783000000001,0,20.25,0,0,None,1500,0,0,0,0,53,0,0.0,1508.38,0.0,1048.45,1,0,92561
3818,0,0,1,0,58,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),109.1,6393.65,0,51,7,37.15,4935,0,Murrieta,0,0,Fiber Optic,33.548869,-117.33416499999998,1,109.1,0,6,None,36149,1,0,1,1,58,2,448.0,2154.7,0.0,6393.65,0,0,92562
3819,1,0,0,0,46,0,No phone service,DSL,1,0,0,0,One year,1,Bank transfer (automatic),30.75,1489.3,0,44,19,0.0,5646,0,Murrieta,0,1,Fiber Optic,33.581045,-117.14719,0,30.75,0,0,None,18311,0,0,0,0,46,0,0.0,0.0,0.0,1489.3,0,1,92563
3820,1,1,1,0,72,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),112.9,8061.5,0,69,14,30.3,5569,0,Nuevo,1,1,Cable,33.827690000000004,-117.102244,1,112.9,0,6,Offer A,7344,1,0,1,1,72,3,1129.0,2181.6,0.0,8061.5,0,0,92567
3821,0,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.2,74.2,1,70,25,48.95,4684,1,Perris,0,0,Cable,33.787298,-117.320676,0,77.168,0,0,Offer E,36817,0,1,0,0,1,6,0.0,48.95,0.0,74.2,0,0,92570
3822,0,0,1,1,6,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Mailed check,94.05,518.75,0,39,19,41.29,3083,0,Perris,1,0,Fiber Optic,33.828289,-117.20166599999999,1,94.05,2,7,None,26357,0,0,1,0,6,4,99.0,247.74,0.0,518.75,0,0,92571
3823,1,0,1,0,72,1,1,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),78.85,5763.15,0,24,85,39.61,5091,0,San Jacinto,1,1,Fiber Optic,33.806708,-117.02006999999999,1,78.85,0,2,Offer A,4456,1,0,1,1,72,2,4899.0,2851.92,0.0,5763.15,1,0,92582
3824,1,0,0,0,4,1,0,DSL,0,0,0,1,Month-to-month,1,Mailed check,55.3,238.5,0,33,3,21.03,3684,0,San Jacinto,0,1,Fiber Optic,33.796568,-116.924723,0,55.3,0,0,None,21349,0,0,0,1,4,0,0.72,84.12,0.0,238.5,0,1,92583
3825,0,0,1,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.35,1031.7,0,44,0,9.87,5699,0,Menifee,0,0,NA,33.653338,-117.178271,1,19.35,2,3,None,14068,0,0,1,0,52,0,0.0,513.24,0.0,1031.7,0,0,92584
3826,1,0,1,1,0,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.35, ,0,22,0,36.37,2299,0,Sun City,0,1,NA,33.739412,-117.17333400000001,1,25.35,2,3,None,8692,0,2,1,0,10,2,0.0,363.7,0.0,253.5,1,0,92585
3827,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.45,34.8,0,23,0,46.0,4196,0,Sun City,0,0,NA,33.707483,-117.200006,0,20.45,0,0,None,18161,0,0,0,0,2,0,0.0,92.0,0.0,34.8,1,0,92586
3828,0,0,1,0,65,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.35,1319.95,0,29,0,48.66,5076,0,Sun City,0,0,NA,33.69887,-117.25071000000001,1,19.35,0,7,Offer B,13151,0,0,1,0,65,1,0.0,3162.9,0.0,1319.95,1,0,92587
3829,1,1,1,0,43,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.0,4388.4,1,68,22,31.25,3123,1,Temecula,0,1,DSL,33.475493,-117.219551,1,105.04,0,8,Offer B,3070,0,1,1,0,43,4,0.0,1343.75,0.0,4388.4,0,1,92590
3830,1,0,1,0,4,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.2,420.2,1,57,11,28.22,2650,1,Temecula,0,1,Fiber Optic,33.540603999999995,-117.10909,1,104.208,0,1,None,25655,0,1,1,1,4,8,46.0,112.88,0.0,420.2,0,0,92591
3831,1,1,1,0,25,1,1,Fiber optic,1,0,0,1,One year,1,Electronic check,89.05,2177.45,1,80,28,33.63,2673,1,Temecula,0,1,Cable,33.507255,-117.029473,1,92.61200000000001,0,3,Offer C,46171,0,0,1,0,25,6,610.0,840.7500000000001,0.0,2177.45,0,0,92592
3832,0,0,1,0,51,1,1,DSL,0,1,1,1,One year,1,Credit card (automatic),78.65,3950.85,0,35,4,25.45,5408,0,Wildomar,0,0,DSL,33.617108,-117.253349,1,78.65,0,10,Offer B,19368,1,0,1,1,51,0,15.8,1297.95,0.0,3950.85,0,1,92595
3833,1,0,0,0,12,1,1,DSL,0,0,1,1,Month-to-month,0,Bank transfer (automatic),74.75,827.05,0,21,53,18.52,3521,0,Winchester,1,1,DSL,33.657433000000005,-117.04253999999999,0,74.75,0,0,None,4093,0,0,0,1,12,0,0.0,222.24,0.0,827.05,1,1,92596
3834,0,0,1,1,57,1,0,DSL,1,0,1,1,One year,1,Bank transfer (automatic),70.1,3913.3,1,46,8,36.65,4669,1,Irvine,0,0,Cable,33.720359,-117.733655,1,72.904,0,1,Offer B,2762,0,2,1,1,57,1,313.0,2089.05,0.0,3913.3,0,0,92602
3835,0,0,1,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.9,533.5,0,38,0,4.47,4158,0,Irvine,0,0,NA,33.688546,-117.788091,1,19.9,3,1,Offer C,27369,0,0,1,0,24,2,0.0,107.28,0.0,533.5,0,0,92604
3836,0,0,1,0,64,1,1,DSL,0,0,0,0,One year,0,Bank transfer (automatic),58.35,3756.45,0,27,52,40.28,5331,0,Irvine,1,0,Fiber Optic,33.703976000000004,-117.82417199999999,1,58.35,0,1,Offer B,17621,1,0,1,0,64,3,1953.0,2577.92,0.0,3756.45,1,0,92606
3837,0,0,0,0,4,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,105.65,443.9,1,29,57,43.45,4663,1,Foothill Ranch,1,0,Fiber Optic,33.698728,-117.67768000000001,0,109.876,0,0,None,10936,1,0,0,1,4,4,0.0,173.8,0.0,443.9,1,1,92610
3838,0,0,0,0,26,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),100.5,2599.95,0,60,3,25.66,2921,0,Irvine,1,0,Fiber Optic,33.643095,-117.810896,0,100.5,0,0,Offer C,41062,0,0,0,1,26,1,0.0,667.16,0.0,2599.95,0,1,92612
3839,0,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,284.3,0,57,0,37.9,3591,0,Irvine,0,0,NA,33.680302000000005,-117.83329599999999,1,20.05,1,3,None,22499,0,1,1,0,15,1,0.0,568.5,0.0,284.3,0,0,92614
3840,1,1,1,0,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.65,1740.8,0,76,0,29.43,6469,0,Irvine,0,1,NA,33.667145,-117.73213500000001,1,25.65,0,0,None,6301,0,0,0,0,64,0,0.0,1883.52,0.0,1740.8,0,0,92618
3841,1,1,1,0,36,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,96.5,3436.1,1,77,3,16.61,4652,1,Irvine,0,1,DSL,33.716136,-117.752574,1,100.36,0,1,None,26419,0,0,1,0,36,3,0.0,597.96,0.0,3436.1,0,1,92620
3842,0,0,1,0,27,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Credit card (automatic),95.0,2462.55,0,21,26,18.42,4235,0,Capistrano Beach,0,0,Fiber Optic,33.458754,-117.665104,1,95.0,0,1,Offer C,7465,0,0,1,1,27,1,640.0,497.34,0.0,2462.55,1,0,92624
3843,1,1,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.85,70.85,1,65,14,49.6,3022,1,Corona Del Mar,0,1,DSL,33.600986999999996,-117.862734,1,73.684,0,1,Offer E,13422,0,2,1,0,1,1,0.0,49.6,0.0,70.85,0,0,92625
3844,0,0,0,0,35,1,1,DSL,1,0,1,1,One year,1,Credit card (automatic),85.95,3110.1,1,27,51,8.8,3833,1,Costa Mesa,1,0,Cable,33.678591,-117.90547099999999,0,89.38799999999999,0,0,Offer C,48207,1,0,0,1,35,4,1586.0,308.0,0.0,3110.1,1,0,92626
3845,1,0,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.9,280.85,1,50,33,33.65,4479,1,Costa Mesa,1,1,Cable,33.645672,-117.92261299999998,0,76.85600000000002,0,0,Offer E,62069,0,1,0,0,4,2,0.0,134.6,0.0,280.85,0,1,92627
3846,0,0,1,1,8,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.45,411.75,0,30,51,5.09,4651,0,Dana Point,0,0,Cable,33.477923,-117.70531399999999,1,45.45,2,0,Offer E,27730,0,1,0,0,8,2,210.0,40.72,0.0,411.75,0,0,92629
3847,1,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.0,198.6,0,51,0,19.1,4802,0,Lake Forest,0,1,NA,33.644849,-117.68425400000001,0,20.0,0,0,Offer D,59176,0,1,0,0,10,1,0.0,191.0,0.0,198.6,0,0,92630
3848,0,0,0,0,2,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,49.2,103.7,0,44,4,29.28,2342,0,Huntington Beach,0,0,DSL,33.666301000000004,-117.969501,0,49.2,0,0,Offer E,56517,0,0,0,0,2,1,0.0,58.56,0.0,103.7,0,1,92646
3849,0,0,1,0,58,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),109.45,6144.55,1,39,26,27.99,6424,1,Huntington Beach,1,0,Fiber Optic,33.723579,-118.00544099999999,1,113.82799999999999,0,1,Offer B,58764,0,2,1,1,58,2,1598.0,1623.4199999999996,0.0,6144.55,0,0,92647
3850,1,0,1,0,51,1,0,DSL,1,1,1,1,Two year,1,Credit card (automatic),83.25,4089.45,0,33,9,40.34,5340,0,Huntington Beach,1,1,DSL,33.679659,-118.016195,1,83.25,0,1,Offer B,42663,1,0,1,1,51,1,0.0,2057.34,0.0,4089.45,0,1,92648
3851,0,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.25,864.2,0,52,0,24.33,5596,0,Huntington Beach,0,0,NA,33.721917,-118.043237,1,19.25,2,1,Offer B,32304,0,0,1,0,46,1,0.0,1119.1799999999996,0.0,864.2,0,0,92649
3852,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.65,19.65,0,40,0,13.85,3075,0,Laguna Beach,0,1,NA,33.570023,-117.773669,0,19.65,0,0,Offer E,25206,0,0,0,0,1,2,0.0,13.85,0.0,19.65,0,0,92651
3853,1,0,0,0,46,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),72.8,3249.4,0,38,26,41.1,2642,0,Laguna Hills,0,1,Fiber Optic,33.606899,-117.717854,0,72.8,0,0,Offer B,48273,0,0,0,0,46,0,845.0,1890.6,0.0,3249.4,0,0,92653
3854,0,0,1,0,50,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),109.65,5405.8,0,62,13,34.57,4676,0,Midway City,0,0,DSL,33.744439,-117.98588000000001,1,109.65,0,4,Offer B,8660,1,0,1,1,50,1,0.0,1728.5,0.0,5405.8,0,1,92655
3855,1,0,1,1,53,1,0,DSL,0,1,1,0,Month-to-month,0,Credit card (automatic),65.0,3363.8,0,31,19,2.11,5534,0,Aliso Viejo,0,1,Fiber Optic,33.571259000000005,-117.731917,1,65.0,1,9,Offer B,41237,1,1,1,0,53,1,639.0,111.83,0.0,3363.8,0,0,92656
3856,1,0,1,0,61,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,114.1,7132.15,0,48,7,12.32,5239,0,Newport Coast,1,1,DSL,33.603282,-117.82184099999999,1,114.1,0,8,Offer B,5597,1,0,1,1,61,0,0.0,751.52,0.0,7132.15,0,1,92657
3857,1,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.65,93.55,0,40,0,42.52,5597,0,Newport Beach,0,1,NA,33.634626000000004,-117.874882,0,20.65,0,0,Offer E,28687,0,0,0,0,5,0,0.0,212.6,0.0,93.55,0,0,92660
3858,1,0,0,0,47,1,0,DSL,1,1,1,1,One year,1,Bank transfer (automatic),86.95,4138.9,0,33,25,36.78,5631,0,Newport Beach,1,1,DSL,33.601309,-117.902304,0,86.95,0,0,Offer B,4242,1,1,0,1,47,1,0.0,1728.66,0.0,4138.9,0,1,92661
3859,0,0,0,0,54,1,1,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),94.75,5121.75,0,30,30,37.65,5665,0,Newport Beach,1,0,Fiber Optic,33.606336,-117.893042,0,94.75,0,0,Offer B,3124,0,0,0,0,54,3,153.65,2033.1,0.0,5121.75,0,1,92662
3860,1,0,0,1,19,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),25.35,566.1,0,19,59,0.0,3072,0,Newport Beach,0,1,DSL,33.62251,-117.927024,0,25.35,2,0,Offer D,22133,0,0,0,1,19,1,0.0,0.0,0.0,566.1,1,1,92663
3861,0,0,0,1,26,1,0,Fiber optic,0,1,1,1,Two year,1,Electronic check,105.45,2715.3,0,63,19,2.48,5980,0,San Clemente,1,0,Fiber Optic,33.429488,-117.60943200000001,0,105.45,1,0,Offer C,34946,1,0,0,1,26,1,0.0,64.48,0.0,2715.3,0,1,92672
3862,1,0,1,1,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.4,1782.05,0,31,0,9.33,4954,0,San Clemente,0,1,NA,33.4725,-117.584273,1,25.4,1,10,Offer A,15297,0,0,1,0,70,2,0.0,653.1,0.0,1782.05,0,0,92673
3863,1,0,1,0,17,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,102.55,1742.5,0,58,2,10.11,3803,0,San Juan Capistrano,1,1,DSL,33.521446999999995,-117.60255500000001,1,102.55,0,2,Offer D,34321,0,0,1,1,17,0,0.0,171.87,0.0,1742.5,0,1,92675
3864,0,0,0,0,30,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.2,2983.8,1,21,90,11.73,3598,1,Silverado,0,0,DSL,33.782346000000004,-117.635263,0,104.208,0,0,Offer C,1859,0,6,0,1,30,3,2685.0,351.9000000000001,0.0,2983.8,1,0,92676
3865,0,0,0,1,1,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,24.0,24,0,45,0,32.95,2559,0,Laguna Niguel,0,0,NA,33.529047,-117.701175,0,24.0,1,0,Offer E,62103,0,0,0,0,1,1,0.0,32.95,0.0,24.0,0,0,92677
3866,0,0,1,1,19,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.6,485.9,0,50,0,38.43,5038,0,Trabuco Canyon,0,0,NA,33.631119,-117.567346,1,25.6,2,4,Offer D,32268,0,0,1,0,19,0,0.0,730.17,0.0,485.9,0,0,92679
3867,0,0,1,0,26,1,0,DSL,0,1,1,1,Two year,1,Credit card (automatic),73.5,1905.7,0,23,58,34.12,3596,0,Westminster,1,0,Fiber Optic,33.752590999999995,-117.99366100000002,1,73.5,0,6,Offer C,88230,0,0,1,1,26,1,1105.0,887.1199999999999,17.03,1905.7,1,0,92683
3868,0,0,1,1,21,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),74.05,1565.7,1,32,29,5.07,5630,1,Rancho Santa Margarita,0,0,DSL,33.624654,-117.611733,1,77.012,0,1,None,42193,0,0,1,0,21,5,454.0,106.47,0.0,1565.7,0,0,92688
3869,1,0,1,0,50,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,98.25,4858.7,0,46,16,38.29,5154,0,Mission Viejo,0,1,Fiber Optic,33.611945,-117.66586699999999,1,98.25,0,10,Offer B,46371,0,0,1,1,50,2,777.0,1914.5,3.55,4858.7,0,0,92691
3870,0,0,1,0,68,0,No phone service,DSL,1,0,1,1,One year,1,Electronic check,54.4,3723.65,0,58,11,0.0,4897,0,Mission Viejo,1,0,DSL,33.60693,-117.644253,1,54.4,0,8,Offer A,46227,0,0,1,1,68,2,410.0,0.0,25.62,3723.65,0,0,92692
3871,1,0,0,0,3,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),101.55,298.35,1,57,7,21.86,4480,1,Ladera Ranch,1,1,Fiber Optic,33.569186,-117.640055,0,105.61200000000001,0,0,Offer E,350,0,3,0,1,3,5,21.0,65.58,0.0,298.35,0,0,92694
3872,1,0,1,1,9,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,103.1,970.45,0,32,57,44.37,4171,0,Santa Ana,1,1,Fiber Optic,33.748478000000006,-117.85891799999999,1,103.1,3,10,Offer E,58157,1,0,1,1,9,3,0.0,399.33,18.62,970.45,0,1,92701
3873,0,0,1,1,51,0,No phone service,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),34.2,1782,0,23,27,0.0,6404,0,Santa Ana,0,0,Cable,33.748635,-117.906125,1,34.2,2,7,Offer B,70011,1,0,1,1,51,0,0.0,0.0,9.39,1782.0,1,1,92703
3874,0,0,0,0,9,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,43.75,405.7,0,48,29,40.73,5644,0,Santa Ana,0,0,DSL,33.719869,-117.907063,0,43.75,0,0,None,91188,0,0,0,0,9,0,118.0,366.57,5.9,405.7,0,0,92704
3875,1,1,1,1,41,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,111.95,4534.9,1,66,32,45.04,3711,1,Santa Ana,1,1,Cable,33.766003999999995,-117.786763,1,116.428,0,1,Offer B,44117,1,0,1,0,41,0,0.0,1846.64,0.0,4534.9,0,1,92705
3876,1,0,0,0,22,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.65,2415.95,0,26,73,28.42,4094,0,Santa Ana,0,1,Fiber Optic,33.765893,-117.881533,0,100.65,0,0,Offer D,37879,0,0,0,1,22,2,0.0,625.24,5.01,2415.95,1,1,92706
3877,0,0,1,1,21,0,No phone service,DSL,1,0,1,1,One year,1,Electronic check,55.95,1157.05,1,30,76,0.0,5531,1,Santa Ana,1,0,Fiber Optic,33.714828999999995,-117.872941,1,58.188,0,1,None,62634,0,0,1,1,21,4,879.0,0.0,0.0,1157.05,0,0,92707
3878,1,0,1,1,71,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),116.05,8297.5,0,41,18,26.38,6481,0,Fountain Valley,1,1,Cable,33.712036,-117.95011299999999,1,116.05,1,5,Offer A,54548,1,0,1,1,71,2,1494.0,1872.98,42.57,8297.5,0,0,92708
3879,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.75,45.75,1,36,31,24.24,3531,1,Tustin,0,1,DSL,33.735802,-117.818805,0,47.58,0,0,None,55062,0,2,0,0,1,5,0.0,24.24,0.0,45.75,0,0,92780
3880,1,0,1,1,26,1,1,DSL,0,0,1,1,One year,1,Credit card (automatic),82.0,2083.1,0,51,57,36.71,3973,0,Tustin,1,1,DSL,33.738543,-117.785046,1,82.0,3,2,Offer C,17494,1,0,1,1,26,0,1187.0,954.46,42.43,2083.1,0,0,92782
3881,1,0,1,0,71,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),65.15,4681.75,0,29,69,40.63,4384,0,Anaheim,0,1,Fiber Optic,33.844983,-117.952151,1,65.15,0,2,Offer A,60553,1,0,1,1,71,1,3230.0,2884.73,4.7,4681.75,1,0,92801
3882,1,0,0,0,4,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),44.8,176.2,0,28,41,43.77,5565,0,Anaheim,0,1,Fiber Optic,33.807864,-117.923782,0,44.8,0,0,Offer E,45086,0,0,0,1,4,2,0.0,175.08,0.0,176.2,1,1,92802
3883,0,0,0,0,12,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,79.8,1001.2,0,61,14,14.42,5906,0,Anaheim,0,0,Fiber Optic,33.818000000000005,-117.974404,0,79.8,0,0,Offer D,81333,0,0,0,0,12,0,140.0,173.04,21.53,1001.2,0,0,92804
3884,0,0,1,0,18,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,88.85,1594.75,0,23,59,18.55,3127,0,Anaheim,0,0,Cable,33.830209,-117.906099,1,88.85,0,8,Offer D,68802,1,0,1,1,18,1,94.09,333.9000000000001,21.58,1594.75,1,1,92805
3885,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.95,212.4,0,42,8,1.64,3641,0,Anaheim,0,0,DSL,33.837959999999995,-117.870494,0,74.95,0,0,Offer E,34398,0,1,0,0,3,2,17.0,4.92,27.6,212.4,0,0,92806
3886,0,1,1,0,72,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),106.85,7677.4,0,69,20,7.85,4768,0,Anaheim,0,0,Fiber Optic,33.848733,-117.788357,1,106.85,0,8,Offer A,36301,0,0,1,1,72,1,153.55,565.1999999999998,0.0,7677.4,0,1,92807
3887,1,0,0,0,11,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,74.95,815.5,1,41,32,25.24,4251,1,Anaheim,0,1,Cable,33.850452000000004,-117.72666799999999,0,77.94800000000002,0,0,None,19629,0,2,0,0,11,3,261.0,277.64,0.0,815.5,0,0,92808
3888,0,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Credit card (automatic),80.15,80.15,1,53,12,4.67,3947,1,Brea,0,0,Cable,33.930199,-117.862898,0,83.35600000000002,0,0,Offer E,34055,0,1,0,1,1,3,0.0,4.67,0.0,80.15,0,1,92821
3889,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.3,259.65,0,44,0,45.03,2823,0,Brea,0,1,NA,33.924143,-117.79387,0,19.3,0,0,Offer D,1408,0,0,0,0,13,2,0.0,585.39,35.28,259.65,0,0,92823
3890,0,0,1,0,72,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,109.25,8109.8,1,57,12,31.13,4261,1,Fullerton,1,0,DSL,33.879983,-117.895482,1,113.62,0,1,None,34592,1,3,1,1,72,3,973.0,2241.36,0.0,8109.8,0,0,92831
3891,1,0,1,0,42,1,1,DSL,1,0,0,0,One year,0,Credit card (automatic),56.1,2386.85,0,56,25,20.65,5904,0,Fullerton,0,1,Fiber Optic,33.868316,-117.929029,1,56.1,0,1,Offer B,24502,0,0,1,0,42,0,59.67,867.3,28.83,2386.85,0,1,92832
3892,0,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.7,340.35,0,27,0,22.26,4222,0,Fullerton,0,0,NA,33.877639,-117.96121200000002,0,19.7,0,0,Offer D,46105,0,0,0,0,17,1,0.0,378.42,0.0,340.35,1,0,92833
3893,0,1,0,0,7,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,51.3,419.35,0,73,18,11.01,3660,0,Fullerton,0,0,DSL,33.902211,-117.914922,0,51.3,0,0,None,21157,0,0,0,0,7,0,75.0,77.07,0.0,419.35,0,0,92835
3894,0,0,1,0,68,1,1,Fiber optic,1,1,1,1,Two year,0,Mailed check,118.6,7990.05,0,27,27,1.29,4175,0,Garden Grove,1,0,DSL,33.787165,-117.93188899999998,1,118.6,0,1,Offer A,50641,1,0,1,1,68,0,0.0,87.72,38.57,7990.05,1,1,92840
3895,1,0,1,1,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.15,1402.25,0,54,0,37.67,5137,0,Garden Grove,0,1,NA,33.786738,-117.982564,1,24.15,2,1,Offer B,31428,0,0,1,0,56,0,0.0,2109.52,29.41,1402.25,0,0,92841
3896,0,0,1,1,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.3,749.35,0,52,0,44.32,4686,0,Garden Grove,0,0,NA,33.764018,-117.93150700000001,1,20.3,3,1,Offer C,43491,0,0,1,0,38,0,0.0,1684.16,10.65,749.35,0,0,92843
3897,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,115.5,8425.15,0,53,10,36.82,4017,0,Garden Grove,1,0,Fiber Optic,33.766476000000004,-117.96979499999999,1,115.5,1,1,Offer A,23481,1,0,1,1,72,1,0.0,2651.04,42.29,8425.15,0,1,92844
3898,0,0,0,0,48,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),25.05,1171.5,0,44,0,34.96,3642,0,Garden Grove,0,0,NA,33.782955,-118.02645600000001,0,25.05,0,0,Offer B,15878,0,0,0,0,48,0,0.0,1678.08,16.38,1171.5,0,0,92845
3899,0,1,1,0,52,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,109.1,5647.95,0,67,17,4.11,4428,0,Norco,1,0,Cable,33.925833000000004,-117.55963899999999,1,109.1,0,1,None,22443,0,0,1,0,52,0,960.0,213.72000000000003,0.0,5647.95,0,0,92860
3900,0,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.65,708.8,0,30,0,18.29,3739,0,Villa Park,0,0,NA,33.817473,-117.81046200000002,1,19.65,2,1,Offer C,5935,0,0,1,0,35,0,0.0,640.15,0.0,708.8,0,0,92861
3901,1,0,1,0,67,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),111.3,7567.2,0,60,30,21.71,4469,0,Orange,1,1,Fiber Optic,33.828779,-117.848299,1,111.3,0,1,Offer A,18058,1,0,1,1,67,0,0.0,1454.5700000000004,36.66,7567.2,0,1,92865
3902,0,0,0,0,1,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,29.9,29.9,0,42,24,0.0,4155,0,Orange,0,0,Cable,33.784597,-117.84453500000001,0,29.9,0,0,None,15396,0,0,0,0,1,0,0.0,0.0,0.0,29.9,0,1,92866
3903,1,0,0,0,53,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,80.6,4348.1,0,56,29,49.21,6113,0,Orange,0,1,DSL,33.81859,-117.821288,0,80.6,0,0,Offer B,40915,1,0,0,0,53,1,0.0,2608.13,39.45,4348.1,0,1,92867
3904,1,0,1,1,34,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.8,635.9,0,44,0,44.54,4985,0,Orange,0,1,NA,33.787796,-117.875928,1,20.8,1,1,Offer C,23172,0,0,1,0,34,0,0.0,1514.36,46.07,635.9,0,0,92868
3905,0,0,0,0,3,0,No phone service,DSL,0,0,1,0,Month-to-month,0,Credit card (automatic),35.2,108.95,1,20,33,0.0,5450,1,Orange,0,0,DSL,33.792790999999994,-117.789749,0,36.608,0,0,Offer E,37916,0,1,0,0,3,1,0.0,0.0,0.0,108.95,1,1,92869
3906,0,0,1,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,78.8,78.8,1,55,33,28.04,5075,1,Placentia,0,0,Fiber Optic,33.881158,-117.85478300000001,1,81.95200000000001,0,1,Offer E,48170,0,0,1,0,1,0,0.0,28.04,0.0,78.8,0,0,92870
3907,1,0,0,0,19,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Mailed check,89.95,1682.4,0,49,6,9.55,3402,0,Corona,1,1,Fiber Optic,33.893823,-117.531446,0,89.95,0,0,Offer D,44875,1,0,0,0,19,2,101.0,181.45,29.64,1682.4,0,0,92879
3908,0,1,1,0,60,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),116.05,6925.9,0,70,11,4.06,4734,0,Corona,1,0,Cable,33.918043,-117.61780900000001,1,116.05,0,1,None,16998,1,0,1,0,60,2,762.0,243.6,0.0,6925.9,0,0,92880
3909,1,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.55,223.15,0,45,0,17.12,5433,0,Corona,0,1,NA,33.833686,-117.51306299999999,0,19.55,0,0,Offer D,21911,0,0,0,0,11,0,0.0,188.32,26.32,223.15,0,0,92881
3910,0,0,0,0,47,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.4,5127.95,1,42,28,35.97,4804,1,Corona,1,0,Cable,33.819385,-117.60021299999998,0,110.656,0,0,Offer B,60294,0,4,0,1,47,1,1436.0,1690.59,0.0,5127.95,0,0,92882
3911,1,0,0,0,18,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,49.4,874.8,1,31,3,20.86,4028,1,Corona,0,1,DSL,33.762351,-117.488725,0,51.376000000000005,0,0,None,13188,0,0,0,0,18,3,26.0,375.48,0.0,874.8,0,0,92883
3912,0,0,1,1,60,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),115.25,6758.45,0,41,28,43.33,5328,0,Yorba Linda,1,0,DSL,33.897253000000006,-117.792202,1,115.25,1,1,Offer B,39458,1,0,1,1,60,0,0.0,2599.8,11.85,6758.45,0,1,92886
3913,1,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.8,1874.3,0,38,0,13.72,6251,0,Yorba Linda,0,1,NA,33.884073,-117.732197,1,24.8,0,1,None,20893,0,0,1,0,72,0,0.0,987.84,16.26,1874.3,0,0,92887
3914,1,0,0,0,39,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.9,791.15,0,26,0,48.02,4041,0,Ventura,0,1,NA,34.360261,-119.30638300000001,0,19.9,0,0,Offer C,32899,0,0,0,0,39,0,0.0,1872.78,20.17,791.15,1,0,93001
3915,0,0,1,0,59,1,0,Fiber optic,1,0,0,0,One year,1,Credit card (automatic),81.25,4639.45,0,43,12,29.6,4709,0,Ventura,1,0,DSL,34.279221,-119.22143700000001,1,81.25,0,1,None,46894,0,0,1,0,59,0,0.0,1746.4,0.0,4639.45,0,1,93003
3916,1,0,1,1,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,69.95,143.9,0,48,19,29.1,5010,0,Ventura,0,1,Fiber Optic,34.278696999999994,-119.167798,1,69.95,2,6,Offer E,27381,0,0,1,0,2,0,2.73,58.2,0.0,143.9,0,1,93004
3917,1,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.1,69.1,1,70,13,16.19,2767,1,Camarillo,0,1,DSL,34.227846,-119.079903,0,71.86399999999998,0,0,None,42853,0,0,0,0,1,2,0.0,16.19,0.0,69.1,0,1,93010
3918,1,0,1,1,20,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.2,1776.55,1,63,11,49.69,2058,1,Camarillo,0,1,DSL,34.205504,-118.99311100000001,1,93.80799999999999,0,1,None,24945,0,0,1,1,20,0,0.0,993.8,0.0,1776.55,0,1,93012
3919,0,0,0,0,6,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),93.55,536.4,1,42,6,43.8,5617,1,Carpinteria,0,0,Cable,34.441398,-119.51316299999999,0,97.292,0,0,Offer E,17409,0,2,0,1,6,2,32.0,262.79999999999995,0.0,536.4,0,0,93013
3920,1,0,0,0,71,1,1,Fiber optic,0,0,0,0,Two year,1,Credit card (automatic),86.4,6172,0,53,15,6.75,4069,0,Fillmore,1,1,DSL,34.408161,-118.86511100000001,0,86.4,0,0,None,16013,1,0,0,0,71,2,926.0,479.25,0.0,6172.0,0,0,93015
3921,0,0,1,0,24,1,1,DSL,1,1,0,0,Month-to-month,0,Mailed check,66.3,1559.45,0,21,27,9.3,2235,0,Moorpark,1,0,Fiber Optic,34.312945,-118.85816899999999,1,66.3,0,6,None,32984,0,0,1,0,24,1,421.0,223.2,32.59,1559.45,1,0,93021
3922,1,1,1,0,67,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),94.65,6079,0,79,23,7.2,4228,0,Oak View,0,1,DSL,34.404544,-119.302118,1,94.65,0,4,Offer A,6503,0,0,1,0,67,0,0.0,482.4,0.0,6079.0,0,1,93022
3923,1,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Mailed check,80.85,80.85,1,64,23,14.91,3096,1,Ojai,0,1,DSL,34.581308,-118.93194799999999,0,84.084,0,0,None,21633,0,1,0,1,1,3,0.0,14.91,0.0,80.85,0,0,93023
3924,0,0,1,1,48,1,1,Fiber optic,0,0,0,1,One year,1,Mailed check,82.05,4029.95,1,41,33,23.95,3365,1,Oxnard,0,0,Cable,34.223244,-119.18012,1,85.33200000000001,0,1,Offer B,79736,0,0,1,1,48,1,1330.0,1149.6,0.0,4029.95,0,0,93030
3925,0,0,1,0,37,1,1,DSL,0,1,0,1,One year,0,Mailed check,72.1,2658.4,0,41,23,42.45,2703,0,Oxnard,0,0,Fiber Optic,34.156628999999995,-119.117218,1,72.1,0,4,None,77791,1,0,1,1,37,0,0.0,1570.65,16.36,2658.4,0,1,93033
3926,1,0,0,0,11,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Mailed check,34.7,383.55,0,60,22,0.0,4310,0,Oxnard,1,1,Fiber Optic,34.184540000000005,-119.22466599999998,0,34.7,0,0,Offer D,25322,0,1,0,0,11,1,0.0,0.0,22.53,383.55,0,1,93035
3927,1,0,1,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.55,51.15,1,41,0,37.61,4115,1,Piru,0,1,NA,34.432843,-118.730106,1,20.55,0,1,Offer E,1459,0,0,1,0,3,4,0.0,112.83,0.0,51.15,0,0,93040
3928,0,0,1,0,18,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),95.95,1745.5,0,56,7,29.6,5009,0,Port Hueneme,1,0,Fiber Optic,34.110124,-119.100972,1,95.95,0,9,Offer D,25634,0,0,1,1,18,2,12.22,532.8000000000002,6.72,1745.5,0,1,93041
3929,1,0,1,1,50,1,0,DSL,0,0,0,0,One year,1,Bank transfer (automatic),44.8,2230.85,0,22,41,36.61,6115,0,Santa Paula,0,1,Fiber Optic,34.402343,-119.094824,1,44.8,2,10,None,32511,0,1,1,0,50,3,0.0,1830.5,36.22,2230.85,1,1,93060
3930,0,0,1,1,67,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,109.4,7281.6,0,53,19,3.3,4103,0,Simi Valley,1,0,Fiber Optic,34.296813,-118.685703,1,109.4,2,7,None,49027,1,0,1,1,67,0,0.0,221.1,38.34,7281.6,0,1,93063
3931,0,0,1,0,25,1,0,DSL,1,1,0,1,Month-to-month,1,Mailed check,71.05,1837.7,0,25,73,2.34,5620,0,Simi Valley,0,0,Fiber Optic,34.269449,-118.76847099999999,1,71.05,0,10,None,64802,1,0,1,1,25,1,0.0,58.5,28.08,1837.7,1,1,93065
3932,0,1,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,78.55,149.55,1,69,15,43.96,5203,1,Somis,1,0,Cable,34.297628,-119.014627,0,81.692,0,0,Offer E,2966,0,0,0,0,2,0,22.0,87.92,0.0,149.55,0,0,93066
3933,1,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.7,180.7,0,37,0,24.89,4194,0,Summerland,0,1,NA,34.420998,-119.60136999999999,0,19.7,0,0,Offer E,576,0,0,0,0,9,3,0.0,224.01,0.0,180.7,0,0,93067
3934,0,0,0,1,10,0,No phone service,DSL,1,1,0,0,One year,0,Mailed check,40.25,411.45,0,52,57,0.0,2876,0,Santa Barbara,0,0,DSL,34.419203,-119.710008,0,40.25,5,0,Offer D,31727,1,0,0,0,10,3,0.0,0.0,17.96,411.45,0,1,93101
3935,0,0,1,0,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.85,1328.35,0,34,0,40.91,4311,0,Santa Barbara,0,0,NA,34.438581,-119.685368,1,19.85,0,0,None,20893,0,0,0,0,70,0,0.0,2863.7,33.29,1328.35,0,0,93103
3936,1,0,0,0,9,1,0,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),68.25,576.95,0,45,24,32.31,4366,0,Santa Barbara,1,1,Cable,34.037341999999995,-119.80078999999999,0,68.25,0,0,Offer E,25771,1,0,0,1,9,0,138.0,290.79,0.0,576.95,0,0,93105
3937,0,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.15,68.45,0,53,0,1.3,5221,0,Santa Barbara,0,0,NA,34.457541,-119.631072,0,20.15,0,0,Offer E,12741,0,0,0,0,4,0,0.0,5.2,0.0,68.45,0,0,93108
3938,0,0,0,0,2,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,50.95,123.05,0,42,24,36.96,5968,0,Santa Barbara,0,0,Fiber Optic,34.406256,-119.72693600000001,0,50.95,0,0,Offer E,10986,0,0,0,0,2,0,0.0,73.92,0.0,123.05,0,1,93109
3939,0,0,0,1,1,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,78.65,78.65,1,41,11,46.09,2728,1,Santa Barbara,0,0,Fiber Optic,34.437945,-119.77191,0,81.796,0,0,Offer E,15757,0,4,0,1,1,2,0.0,46.09,0.0,78.65,0,0,93110
3940,1,0,0,0,19,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),25.15,468.35,0,37,6,0.0,3784,0,Santa Barbara,0,1,Cable,34.460196999999994,-119.80260200000001,0,25.15,0,0,Offer D,16477,0,0,0,0,19,0,0.0,0.0,0.0,468.35,0,1,93111
3941,1,0,1,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.25,174.7,0,22,0,49.83,3149,0,Goleta,0,1,NA,34.489983,-120.091246,1,20.25,3,0,Offer E,49975,0,0,0,0,7,2,0.0,348.81,0.0,174.7,1,0,93117
3942,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,42.9,42.9,1,47,12,4.02,4895,1,Alpaugh,0,1,DSL,35.869626000000004,-119.49877099999999,0,44.61600000000001,0,0,Offer E,1054,0,3,0,0,1,1,0.0,4.02,0.0,42.9,0,0,93201
3943,1,1,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.0,44,0,69,4,28.67,4320,0,Armona,0,1,Fiber Optic,36.315979,-119.710852,0,44.0,0,0,Offer E,2872,0,0,0,0,1,0,0.0,28.67,0.0,44.0,0,1,93202
3944,0,0,1,1,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.25,172.35,0,59,0,12.55,4272,0,Arvin,0,0,NA,35.116307,-118.817644,1,20.25,3,10,None,16206,0,2,1,0,9,1,0.0,112.95,0.0,172.35,0,0,93203
3945,0,0,0,0,3,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,34.25,139.35,1,26,57,0.0,2802,1,Avenal,0,0,DSL,35.916942999999996,-120.129921,0,35.62000000000001,0,0,Offer E,14697,1,0,0,0,3,3,79.0,0.0,0.0,139.35,1,0,93204
3946,0,0,0,0,9,0,No phone service,DSL,1,0,1,1,Month-to-month,0,Mailed check,58.5,539.85,1,30,53,0.0,3032,1,Bodfish,1,0,Cable,35.523990999999995,-118.40043200000001,0,60.84,0,0,Offer E,1954,1,0,0,1,9,1,286.0,0.0,0.0,539.85,0,0,93205
3947,0,0,0,0,5,1,0,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),55.8,300.4,0,42,26,24.83,5104,0,Buttonwillow,1,0,Fiber Optic,35.451402,-119.488413,0,55.8,0,0,None,2078,0,0,0,0,5,1,78.0,124.15,0.0,300.4,0,0,93206
3948,0,0,1,1,56,1,0,Fiber optic,0,0,1,1,One year,0,Bank transfer (automatic),88.9,4968,0,49,28,12.97,4170,0,California Hot Springs,0,0,Fiber Optic,35.865795,-118.69758999999999,1,88.9,1,4,None,226,0,0,1,1,56,0,0.0,726.32,0.0,4968.0,0,1,93207
3949,0,0,0,1,18,1,1,DSL,1,0,0,0,Month-to-month,0,Mailed check,57.65,992.7,0,25,30,17.51,3425,0,Camp Nelson,0,0,DSL,36.057458000000004,-118.591951,0,57.65,2,0,Offer D,191,0,0,0,0,18,2,0.0,315.18,0.0,992.7,1,1,93208
3950,1,1,0,0,49,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.2,4718.25,1,66,2,32.36,5904,1,Coalinga,0,1,Cable,36.186867,-120.38779299999999,0,100.04799999999999,0,0,Offer B,18036,0,0,0,0,49,5,94.0,1585.64,0.0,4718.25,0,0,93210
3951,1,0,1,0,70,1,1,DSL,1,1,1,0,Two year,0,Mailed check,79.15,5536.5,0,40,2,39.35,4408,0,Corcoran,1,1,Fiber Optic,36.04533,-119.532424,1,79.15,0,1,None,23506,1,0,1,0,70,0,0.0,2754.5,0.0,5536.5,0,1,93212
3952,0,0,0,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),108.05,7806.6,0,19,82,10.05,5430,0,Delano,1,0,DSL,35.772244,-119.20968899999998,0,108.05,0,0,None,37280,1,0,0,1,72,3,0.0,723.6,0.0,7806.6,1,1,93215
3953,0,1,0,0,6,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,74.4,434.1,1,75,30,8.91,3964,1,Ducor,1,0,Cable,35.846067,-119.00407299999999,0,77.376,0,0,Offer E,823,0,2,0,0,6,3,130.0,53.46,0.0,434.1,0,0,93218
3954,1,1,1,0,17,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.8,1563.9,0,79,13,46.44,4831,0,Earlimart,0,1,Fiber Optic,35.858053999999996,-119.305858,1,94.8,0,7,None,9318,0,0,1,0,17,2,203.0,789.48,0.0,1563.9,0,0,93219
3955,1,0,1,0,29,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,45.9,1332.4,0,43,15,0.0,5074,0,Exeter,0,1,Fiber Optic,36.301689,-119.01823300000001,1,45.9,0,3,None,13333,0,0,1,1,29,0,19.99,0.0,0.0,1332.4,0,1,93221
3956,0,0,1,0,6,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.3,545.2,1,23,64,27.44,4163,1,Frazier Park,1,0,Fiber Optic,34.907911,-119.23428100000001,1,109.512,0,1,Offer E,1526,0,0,1,1,6,6,349.0,164.64,0.0,545.2,1,0,93222
3957,1,0,1,0,63,1,1,Fiber optic,0,0,1,1,Two year,0,Electronic check,102.6,6296.75,0,35,22,2.72,4004,0,Farmersville,1,1,Cable,36.29878,-119.20102800000001,1,102.6,0,4,None,8644,0,0,1,1,63,1,1385.0,171.36,0.0,6296.75,0,0,93223
3958,1,0,1,0,16,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),73.85,1284.2,1,32,33,17.96,3226,1,Fellows,0,1,Cable,35.215731,-119.57013,1,76.804,0,1,None,626,0,0,1,0,16,2,0.0,287.36,0.0,1284.2,0,1,93224
3959,1,0,0,0,59,1,0,DSL,0,0,0,1,One year,1,Bank transfer (automatic),61.35,3645.5,0,46,6,9.7,6250,0,Frazier Park,1,1,DSL,34.827662,-118.999073,0,61.35,0,0,None,4498,0,0,0,1,59,0,0.0,572.3,0.0,3645.5,0,1,93225
3960,0,0,0,0,3,1,0,DSL,0,0,1,0,Month-to-month,0,Electronic check,57.55,161.45,0,21,42,48.3,4099,0,Glennville,1,0,Cable,35.735694,-118.738483,0,57.55,0,0,None,296,0,0,0,0,3,0,0.0,144.89999999999995,0.0,161.45,1,1,93226
3961,0,0,0,0,8,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Mailed check,29.25,226.95,0,57,2,0.0,2038,0,Hanford,0,0,Fiber Optic,36.292229999999996,-119.622676,0,29.25,0,0,None,53204,0,0,0,0,8,2,0.0,0.0,0.0,226.95,0,1,93230
3962,0,1,1,0,7,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.55,646.85,1,75,13,21.43,5245,1,Huron,0,0,Fiber Optic,36.217864,-120.08011699999999,1,87.932,0,1,Offer E,6918,0,0,1,0,7,4,0.0,150.01,0.0,646.85,0,1,93234
3963,0,0,0,0,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.6,1441.65,0,37,0,32.99,6161,0,Ivanhoe,0,0,NA,36.385818,-119.22424299999999,0,19.6,0,0,None,4517,0,0,0,0,68,1,0.0,2243.32,0.0,1441.65,0,0,93235
3964,0,0,1,1,68,1,1,Fiber optic,1,0,1,1,Two year,0,Credit card (automatic),111.75,7511.3,0,40,57,14.11,4967,0,Kernville,1,0,DSL,35.852892,-118.397782,1,111.75,3,3,None,1873,1,0,1,1,68,0,428.14,959.48,0.0,7511.3,0,1,93238
3965,0,1,1,0,52,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,106.5,5621.85,0,70,18,27.74,4499,0,Kettleman City,1,0,Fiber Optic,35.996922999999995,-120.000951,1,106.5,0,9,None,1809,0,0,1,0,52,0,0.0,1442.48,0.0,5621.85,0,1,93239
3966,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),107.7,7919.8,0,29,85,41.94,4351,0,Lake Isabella,0,1,DSL,35.607875,-118.46631799999999,1,107.7,1,4,None,5564,1,0,1,1,72,2,673.18,3019.68,0.0,7919.8,1,1,93240
3967,0,0,1,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.3,593.2,0,42,0,45.26,5817,0,Lamont,0,0,NA,35.245034999999994,-118.905553,1,19.3,0,1,None,15364,0,0,1,0,32,0,0.0,1448.32,0.0,593.2,0,0,93241
3968,0,0,1,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.05,1423.65,0,44,0,47.24,4747,0,Laton,0,0,NA,36.444232,-119.71828500000001,1,20.05,0,1,None,2900,0,1,1,0,72,2,0.0,3401.28,0.0,1423.65,0,0,93242
3969,1,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),69.95,69.95,0,46,14,11.45,5133,0,Lebec,0,1,Fiber Optic,34.845861,-118.88516299999999,1,69.95,1,10,None,1247,0,0,1,0,1,0,0.0,11.45,0.0,69.95,0,1,93243
3970,1,0,1,1,42,1,0,DSL,1,0,0,1,One year,0,Credit card (automatic),63.7,2763.35,0,29,69,44.95,3764,0,Lemon Cove,0,1,Fiber Optic,36.462671,-118.99729099999999,1,63.7,3,10,None,293,1,0,1,1,42,0,1907.0,1887.9,0.0,2763.35,1,0,93244
3971,0,0,0,0,25,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.75,692.1,1,61,0,19.75,4931,1,Lemoore,0,0,NA,36.303666,-119.825657,0,24.75,0,0,Offer C,30419,0,0,0,0,25,1,0.0,493.75,0.0,692.1,0,0,93245
3972,1,0,0,0,45,1,0,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),50.9,2298.55,0,45,16,19.39,5274,0,Lindsay,0,1,Fiber Optic,36.205465000000004,-119.085807,0,50.9,0,0,None,15508,0,0,0,0,45,2,368.0,872.5500000000002,0.0,2298.55,0,0,93247
3973,0,0,1,1,43,0,No phone service,DSL,1,0,1,1,One year,1,Credit card (automatic),60.4,2640.55,0,46,10,0.0,2725,0,Lost Hills,1,0,Cable,35.637715,-119.893068,1,60.4,2,8,None,2502,1,0,1,1,43,2,0.0,0.0,0.0,2640.55,0,1,93249
3974,1,0,1,0,37,1,1,DSL,1,0,1,1,One year,0,Mailed check,79.25,2911.8,0,43,28,9.26,2322,0,Mc Farland,1,1,Fiber Optic,35.666886,-119.18671699999999,1,79.25,0,6,None,10781,0,0,1,1,37,1,815.0,342.62,0.0,2911.8,0,0,93250
3975,0,1,0,0,20,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),85.8,1727.5,1,67,16,29.29,3336,1,Mc Kittrick,0,0,DSL,35.38381,-119.73088500000001,0,89.23200000000001,0,0,Offer D,302,0,0,0,1,20,1,276.0,585.8,0.0,1727.5,0,0,93251
3976,0,0,0,0,4,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.45,86.6,1,31,10,0.0,4909,1,Temecula,0,0,Cable,33.507255,-117.029473,0,25.428,0,0,Offer E,46171,0,0,0,0,4,3,0.0,0.0,0.0,86.6,0,1,92592
3977,1,0,1,0,63,1,0,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),110.1,6705.7,0,46,15,3.18,6216,0,New Cuyama,1,1,Fiber Optic,34.956577,-119.750142,1,110.1,0,8,None,798,1,0,1,1,63,0,0.0,200.34,0.0,6705.7,0,1,93254
3978,1,0,0,0,3,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Mailed check,90.7,237.65,0,47,10,5.39,3953,0,Temecula,0,1,Fiber Optic,33.507255,-117.029473,0,90.7,0,0,None,46171,0,0,0,1,3,0,0.0,16.169999999999998,0.0,237.65,0,1,92592
3979,1,0,1,1,66,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.3,1672.35,0,59,0,38.55,5617,0,Pixley,0,1,NA,35.957019,-119.330928,1,25.3,3,5,None,4198,0,0,1,0,66,0,0.0,2544.3,0.0,1672.35,0,0,93256
3980,1,0,0,0,28,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.7,2979.5,1,33,14,30.48,2464,1,Porterville,1,1,DSL,36.008958,-118.891593,0,109.928,0,0,Offer C,65566,0,0,0,1,28,0,0.0,853.44,0.0,2979.5,0,1,93257
3981,0,1,0,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,85.2,695.75,0,70,29,44.63,2565,0,Posey,0,0,Fiber Optic,35.861928000000006,-118.636698,0,85.2,0,0,Offer E,266,0,0,0,0,8,0,0.0,357.04,0.0,695.75,0,1,93260
3982,1,0,0,1,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.35,1654.6,0,36,0,4.89,4155,0,Richgrove,0,1,NA,35.809921,-119.12743700000001,0,24.35,3,0,None,2956,0,0,0,0,71,2,0.0,347.19,0.0,1654.6,0,0,93261
3983,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.25,24.25,1,64,8,0.0,2846,1,Sequoia National Park,0,1,Cable,36.527243,-118.59493799999998,0,25.22,0,0,Offer E,56,0,2,0,0,1,3,0.0,0.0,0.0,24.25,0,0,93262
3984,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.1,1857.85,0,43,0,35.62,5611,0,Shafter,0,0,NA,35.490705,-119.286833,1,25.1,2,4,None,15177,0,1,1,0,72,1,0.0,2564.64,0.0,1857.85,0,0,93263
3985,1,1,1,0,16,1,0,DSL,1,1,0,0,Month-to-month,1,Bank transfer (automatic),54.55,825.1,0,79,23,35.53,3324,0,Springville,0,1,DSL,36.245926000000004,-118.69313799999999,1,54.55,0,5,None,3546,0,0,1,0,16,2,190.0,568.48,0.0,825.1,0,0,93265
3986,1,0,1,0,66,1,1,Fiber optic,1,1,0,0,Two year,0,Mailed check,96.6,6424.25,0,43,20,36.55,4454,0,Stratford,1,1,Cable,36.175255,-119.813805,1,96.6,0,5,None,1729,1,0,1,0,66,2,0.0,2412.3,0.0,6424.25,0,1,93266
3987,0,0,0,0,11,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.5,837.95,1,48,4,15.6,2291,1,Strathmore,0,0,DSL,36.141319,-119.129075,0,79.56,0,0,None,5689,0,3,0,0,11,3,34.0,171.6,0.0,837.95,0,0,93267
3988,1,0,0,0,51,1,1,DSL,1,1,1,0,One year,1,Credit card (automatic),81.15,4126.2,0,22,59,34.75,4549,0,Taft,1,1,Fiber Optic,35.184837,-119.402525,0,81.15,0,0,None,14937,1,0,0,0,51,1,243.45,1772.25,0.0,4126.2,1,1,93268
3989,0,0,0,1,8,0,No phone service,DSL,1,0,0,1,Month-to-month,1,Electronic check,38.5,330.8,0,22,51,0.0,4194,0,Terra Bella,0,0,Fiber Optic,35.939068,-119.04366599999999,0,38.5,1,0,None,5868,0,0,0,1,8,0,169.0,0.0,0.0,330.8,1,0,93270
3990,1,0,0,0,14,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,92.9,1337.45,0,47,17,27.8,4296,0,Three Rivers,0,1,Fiber Optic,36.413433000000005,-118.854708,0,92.9,0,0,Offer D,2318,0,0,0,1,14,0,0.0,389.2,0.0,1337.45,0,1,93271
3991,0,0,0,0,4,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,93.5,362.2,1,47,4,7.39,4554,1,Temecula,0,0,DSL,33.507255,-117.029473,0,97.24,0,0,Offer E,46171,1,0,0,1,4,4,0.0,29.56,0.0,362.2,0,1,92592
3992,0,0,0,0,70,1,1,DSL,1,1,1,1,Two year,0,Mailed check,84.7,5991.05,0,44,10,16.93,4180,0,Tulare,1,0,DSL,36.185471,-119.375243,0,84.7,0,0,None,56101,0,0,0,1,70,0,0.0,1185.1,0.0,5991.05,0,1,93274
3993,0,0,0,1,70,1,1,DSL,1,1,0,0,Two year,0,Electronic check,66.0,4891.5,0,54,57,16.75,5265,0,Tupman,0,0,Cable,35.316263,-119.40255900000001,0,66.0,3,0,None,236,1,0,0,0,70,2,2788.0,1172.5,0.0,4891.5,0,0,93276
3994,0,1,1,0,54,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),101.5,5373.1,1,75,9,33.49,6405,1,Visalia,0,0,DSL,36.303793,-119.375646,1,105.56,0,0,Offer B,44741,0,0,0,1,54,1,484.0,1808.46,0.0,5373.1,0,0,93277
3995,1,0,0,1,28,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),74.9,2068.55,1,60,6,44.28,5392,1,Wasco,0,1,Cable,35.652242,-119.4464,0,77.89600000000002,0,0,Offer C,22760,0,0,0,0,28,2,124.0,1239.84,0.0,2068.55,0,0,93280
3996,1,0,0,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.75,487.05,0,40,0,47.51,4117,0,Weldon,0,1,NA,35.556470000000004,-118.244914,0,20.75,0,0,None,1935,0,0,0,0,24,2,0.0,1140.24,0.0,487.05,0,0,93283
3997,0,0,1,0,69,1,0,DSL,0,1,0,1,Two year,1,Credit card (automatic),61.45,4131.2,0,27,69,2.73,4162,0,Wofford Heights,0,0,DSL,35.690535,-118.552784,1,61.45,0,1,None,2515,0,0,1,1,69,3,2851.0,188.37,0.0,4131.2,1,0,93285
3998,1,0,1,1,42,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,54.5,2301.15,0,30,73,18.93,3449,0,Woodlake,0,1,Fiber Optic,36.464634999999994,-119.094348,1,54.5,1,7,None,8870,0,0,1,0,42,1,1680.0,795.06,0.0,2301.15,0,0,93286
3999,0,1,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.6,131.65,1,74,23,15.32,4596,1,Woody,0,0,DSL,35.710244,-118.881679,0,72.384,0,0,Offer E,88,0,1,0,0,2,1,3.03,30.64,0.0,131.65,0,1,93287
4000,0,1,0,0,39,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.75,4036,0,72,13,10.03,3860,0,Visalia,1,0,Fiber Optic,36.391777000000005,-119.37284199999999,0,99.75,0,0,None,36718,0,1,0,0,39,2,52.47,391.17,0.0,4036.0,0,1,93291
4001,1,0,1,1,45,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),109.75,4900.65,0,62,27,7.48,4221,0,Visalia,1,1,DSL,36.37559,-119.21168899999999,1,109.75,3,2,None,30395,1,0,1,1,45,0,1323.0,336.6,0.0,4900.65,0,0,93292
4002,1,0,1,1,72,1,1,DSL,1,1,1,0,Two year,1,Bank transfer (automatic),80.85,5727.45,0,55,12,9.3,6067,0,Bakersfield,1,1,Fiber Optic,35.383937,-119.02042800000001,1,80.85,2,6,None,12963,1,0,1,0,72,0,0.0,669.6,0.0,5727.45,0,1,93301
4003,0,0,0,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.3,743.05,0,43,0,43.19,5919,0,Bakersfield,0,0,NA,35.339796,-119.023552,0,20.3,0,0,None,44588,0,0,0,0,38,1,0.0,1641.2199999999998,0.0,743.05,0,0,93304
4004,1,0,1,0,72,1,1,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),67.8,4804.65,0,46,6,15.52,5242,0,Bakersfield,1,1,Fiber Optic,35.391733,-118.984109,1,67.8,0,1,None,35643,1,0,1,0,72,1,28.83,1117.44,0.0,4804.65,0,1,93305
4005,1,0,0,0,1,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,24.05,24.05,1,21,0,20.26,3162,1,Bakersfield,0,1,NA,35.449881,-118.84144199999999,0,24.05,0,0,None,53481,0,0,0,0,1,2,0.0,20.26,0.0,24.05,1,0,93306
4006,1,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.8,1414.65,0,54,0,38.84,5027,0,Bakersfield,0,1,NA,35.280113,-118.962329,1,19.8,2,10,None,59195,0,0,1,0,72,1,0.0,2796.4800000000005,0.0,1414.65,0,0,93307
4007,1,0,1,0,55,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.7,1443.65,0,54,0,12.21,6228,0,Bakersfield,0,1,NA,35.559616999999996,-118.92518500000001,1,25.7,0,1,None,44915,0,0,1,0,55,2,0.0,671.5500000000002,0.0,1443.65,0,0,93308
4008,0,0,1,1,51,0,No phone service,DSL,0,0,1,1,One year,1,Electronic check,56.15,2898.95,0,42,76,0.0,4132,0,Bakersfield,1,0,Fiber Optic,35.342890999999995,-119.064803,1,56.15,3,4,None,58632,1,0,1,1,51,3,0.0,0.0,0.0,2898.95,0,1,93309
4009,1,0,0,0,63,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),86.7,5309.5,0,24,47,29.58,5841,0,Bakersfield,1,1,Cable,35.16207,-119.19448799999999,0,86.7,0,0,None,20440,1,0,0,1,63,2,2495.0,1863.54,0.0,5309.5,1,0,93311
4010,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,20.4,0,29,0,45.91,2152,0,Bakersfield,0,0,NA,35.392599,-119.245341,0,20.4,0,0,None,40836,0,0,0,0,1,0,0.0,45.91,0.0,20.4,1,0,93312
4011,0,0,1,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.65,451.55,0,24,0,1.88,4896,0,Bakersfield,0,0,NA,35.140938,-119.051348,1,19.65,3,9,Offer D,25126,0,0,1,0,23,0,0.0,43.24,0.0,451.55,1,0,93313
4012,0,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,50.55,50.55,1,36,6,30.96,3420,1,San Luis Obispo,0,0,DSL,35.233745,-120.626442,0,52.572,0,0,None,27047,0,0,0,0,1,0,0.0,30.96,0.0,50.55,0,1,93401
4013,0,0,0,0,2,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,54.35,117.05,0,38,7,25.81,4916,0,Los Osos,0,0,Fiber Optic,35.279984000000006,-120.824288,0,54.35,0,0,None,14859,1,0,0,0,2,2,0.0,51.62,0.0,117.05,0,1,93402
4014,0,1,0,0,52,1,1,Fiber optic,1,1,1,1,Month-to-month,0,Credit card (automatic),108.1,5839.3,0,76,18,11.01,4251,0,San Luis Obispo,1,0,DSL,35.236549,-120.72734399999999,0,108.1,0,0,None,31982,0,0,0,0,52,1,1051.0,572.52,0.0,5839.3,0,0,93405
4015,0,0,0,0,36,1,1,DSL,1,0,0,0,One year,0,Mailed check,54.45,1893.5,0,40,21,25.95,4462,0,Arroyo Grande,0,0,DSL,35.176235999999996,-120.48324299999999,0,54.45,0,0,None,24499,0,0,0,0,36,2,0.0,934.2,0.0,1893.5,0,1,93420
4016,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.35,45.35,0,39,14,12.46,3980,0,Atascadero,0,0,DSL,35.453912,-120.69461000000001,0,45.35,0,0,None,29539,0,0,0,0,1,0,0.0,12.46,0.0,45.35,0,0,93422
4017,0,0,0,0,28,1,1,DSL,1,0,0,0,One year,0,Mailed check,59.0,1654.45,0,35,7,33.05,4891,0,Avila Beach,1,0,Cable,35.186644,-120.728305,0,59.0,0,0,None,812,0,0,0,0,28,0,116.0,925.4,0.0,1654.45,0,0,93424
4018,0,0,1,1,7,1,0,DSL,1,1,1,0,One year,0,Electronic check,69.45,477.05,0,39,29,18.91,3334,0,Bradley,1,0,Fiber Optic,35.842889,-121.00486200000002,1,69.45,3,1,None,1363,0,0,1,0,7,0,0.0,132.37,0.0,477.05,0,1,93426
4019,1,0,0,0,14,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.55,1415.55,1,56,30,36.97,5224,1,Buellton,0,1,Cable,34.631362,-120.23821799999999,0,104.572,0,0,None,4644,0,2,0,1,14,8,425.0,517.5799999999998,0.0,1415.55,0,0,93427
4020,1,1,1,0,72,0,No phone service,DSL,1,1,1,1,Two year,1,Credit card (automatic),64.95,4546,0,70,7,0.0,4049,0,Cambria,1,1,Fiber Optic,35.591387,-121.032256,1,64.95,0,1,Offer A,6526,1,0,1,0,72,1,318.0,0.0,0.0,4546.0,0,0,93428
4021,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.5,20.5,1,47,0,34.57,2398,1,Casmalia,0,0,NA,34.866032000000004,-120.536546,1,20.5,3,0,None,210,0,0,0,0,1,6,0.0,34.57,0.0,20.5,0,0,93429
4022,0,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,18.85,163.2,0,60,0,41.04,5949,0,Cayucos,0,0,NA,35.511833,-120.91871299999998,0,18.85,0,0,Offer D,3220,0,0,0,0,10,0,0.0,410.4,0.0,163.2,0,0,93430
4023,1,0,0,0,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.8,849.9,0,55,0,38.74,3575,0,Creston,0,1,NA,35.480896,-120.469476,0,19.8,0,0,None,1203,0,0,0,0,42,0,0.0,1627.0800000000004,0.0,849.9,0,0,93432
4024,0,0,0,0,7,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),25.05,189.95,0,42,4,0.0,4404,0,Grover Beach,0,0,Fiber Optic,35.120833000000005,-120.61843,0,25.05,0,0,None,13106,0,0,0,0,7,1,8.0,0.0,0.0,189.95,0,0,93433
4025,1,0,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.8,321.9,1,51,32,7.26,5882,1,Guadalupe,1,1,DSL,34.936,-120.594655,0,77.792,0,0,None,5726,0,1,0,0,4,2,0.0,29.04,0.0,321.9,0,1,93434
4026,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),114.3,8058.55,0,43,13,15.94,5879,0,Lompoc,1,1,Fiber Optic,34.601055,-120.38291699999999,1,114.3,1,1,None,51737,1,0,1,1,72,0,0.0,1147.68,0.0,8058.55,0,1,93436
4027,0,0,1,0,20,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.45,482.8,1,44,11,0.0,3298,1,Lompoc,0,0,Cable,34.757477,-120.55050700000001,1,25.428,0,1,None,6165,0,0,1,0,20,2,53.0,0.0,0.0,482.8,0,0,93437
4028,1,0,0,0,63,1,0,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),109.2,7049.75,0,36,17,13.14,4273,0,Los Alamos,1,1,DSL,34.758699,-120.27583899999999,0,109.2,0,0,None,1328,1,0,0,1,63,0,119.85,827.82,0.0,7049.75,0,1,93440
4029,0,0,0,0,56,0,No phone service,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),45.05,2560.1,0,39,19,0.0,5795,0,Los Olivos,1,0,Cable,34.70434,-120.02609,0,45.05,0,0,None,1317,1,0,0,0,56,1,0.0,0.0,0.0,2560.1,0,1,93441
4030,0,0,0,1,5,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,51.0,286.8,0,22,52,40.03,2789,0,Morro Bay,0,0,Fiber Optic,35.369553,-120.76386399999998,0,51.0,1,0,None,10909,1,0,0,0,5,0,149.0,200.15,0.0,286.8,1,0,93442
4031,0,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),110.45,7982.5,0,33,18,46.23,6030,0,Nipomo,1,0,Cable,35.050345,-120.489599,1,110.45,0,1,None,15405,1,0,1,1,72,0,0.0,3328.56,0.0,7982.5,0,1,93444
4032,1,1,1,1,68,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,84.65,5683.6,0,70,13,20.31,6404,0,Oceano,1,1,DSL,35.059695,-120.60474099999999,1,84.65,1,1,Offer A,7435,0,0,1,0,68,0,739.0,1381.08,0.0,5683.6,0,0,93445
4033,1,0,1,1,67,1,0,DSL,1,1,0,0,One year,0,Mailed check,60.05,3994.05,0,43,19,6.53,6148,0,Paso Robles,0,1,DSL,35.634221999999994,-120.72834099999999,1,60.05,2,1,None,35586,1,0,1,0,67,1,0.0,437.51,0.0,3994.05,0,1,93446
4034,1,0,1,1,8,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),44.65,369.15,0,45,75,30.77,5724,0,Pismo Beach,0,1,DSL,35.165668,-120.65584199999999,1,44.65,3,1,None,8564,0,0,1,0,8,0,277.0,246.16,0.0,369.15,0,0,93449
4035,1,0,1,1,52,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),93.25,4631.7,0,49,10,11.3,4740,0,San Ardo,0,1,Fiber Optic,35.996008,-120.85305,1,93.25,1,1,None,670,1,0,1,1,52,0,0.0,587.6,0.0,4631.7,0,1,93450
4036,0,0,1,1,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.25,401.95,0,29,0,35.44,2429,0,San Miguel,0,0,NA,35.886767,-120.60866100000001,1,20.25,1,10,Offer D,2666,0,0,1,0,18,4,0.0,637.92,0.0,401.95,1,0,93451
4037,0,0,1,1,59,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.45,1534.05,0,40,0,42.37,4746,0,San Simeon,0,0,NA,35.746484,-121.223355,1,25.45,2,0,Offer B,471,0,0,0,0,59,2,0.0,2499.83,0.0,1534.05,0,0,93452
4038,0,0,0,0,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.6,1093,0,60,0,47.07,4192,0,Santa Margarita,0,0,NA,35.303926000000004,-120.25656699999999,0,20.6,0,0,Offer B,2687,0,0,0,0,60,0,0.0,2824.2,0.0,1093.0,0,0,93453
4039,1,0,0,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.1,701.3,0,55,6,7.37,5259,0,Santa Maria,0,1,Cable,34.943523,-120.256729,0,94.1,0,0,None,30540,0,0,0,1,7,0,0.0,51.59,0.0,701.3,0,1,93454
4040,1,0,1,1,59,0,No phone service,DSL,1,0,0,0,One year,0,Mailed check,34.8,1980.3,0,59,19,0.0,6300,0,Santa Maria,1,1,Fiber Optic,34.818227,-120.418784,1,34.8,2,0,Offer B,37364,0,0,0,0,59,1,376.0,0.0,0.0,1980.3,0,0,93455
4041,1,0,0,0,46,0,No phone service,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),60.75,2893.4,0,33,13,0.0,2694,0,Santa Maria,1,1,Fiber Optic,34.959340000000005,-120.490081,0,60.75,0,0,Offer B,43684,1,2,0,1,46,1,0.0,0.0,0.0,2893.4,0,1,93458
4042,1,0,0,0,5,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,51.35,262.3,0,39,7,17.16,2893,0,Santa Ynez,0,1,Fiber Optic,34.630356,-120.032564,0,51.35,0,0,Offer E,5710,0,0,0,0,5,2,0.0,85.8,0.0,262.3,0,1,93460
4043,1,1,1,0,59,0,No phone service,DSL,1,0,1,1,Two year,1,Credit card (automatic),64.05,3886.85,0,77,6,0.0,6306,0,Shandon,1,1,Fiber Optic,35.634488,-120.29353400000001,1,64.05,0,3,None,1255,1,0,1,0,59,1,233.0,0.0,0.0,3886.85,0,0,93461
4044,0,0,1,0,70,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),84.8,5917.55,0,53,24,9.28,4032,0,Solvang,1,0,Cable,34.624399,-120.137875,1,84.8,0,7,None,7958,1,0,1,1,70,0,0.0,649.5999999999998,0.0,5917.55,0,1,93463
4045,0,0,0,0,14,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),71.0,914,1,27,57,36.25,3228,1,Templeton,0,0,DSL,35.536115,-120.739231,0,73.84,0,0,None,7918,0,0,0,0,14,1,521.0,507.5,0.0,914.0,1,0,93465
4046,0,0,0,0,44,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.15,2139.1,0,64,22,18.42,5790,0,Mojave,0,0,Fiber Optic,35.097322999999996,-118.17128799999999,0,50.15,0,0,Offer B,4882,0,0,0,0,44,0,471.0,810.48,0.0,2139.1,0,0,93501
4047,0,0,1,0,64,1,1,Fiber optic,1,0,1,0,Two year,1,Credit card (automatic),94.6,5948.7,0,45,13,1.27,5038,0,California City,1,0,Fiber Optic,35.151491,-117.92759699999999,1,94.6,0,7,Offer B,8316,0,0,1,0,64,1,773.0,81.28,0.0,5948.7,0,0,93505
4048,0,0,1,1,58,0,No phone service,DSL,1,0,1,1,Two year,0,Mailed check,59.75,3624.35,0,25,59,0.0,4678,0,Acton,1,0,DSL,34.501452,-118.207862,1,59.75,3,8,Offer B,7831,1,0,1,1,58,1,2138.0,0.0,0.0,3624.35,1,0,93510
4049,0,1,1,0,46,1,1,Fiber optic,0,0,1,1,One year,0,Electronic check,100.25,4753.85,0,71,15,21.46,5453,0,Benton,0,0,DSL,37.653946999999995,-118.231443,1,100.25,0,5,None,340,1,0,1,0,46,0,0.0,987.16,0.0,4753.85,0,1,93512
4050,1,1,1,0,58,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,98.9,5780.7,0,80,4,31.11,4993,0,Big Pine,0,1,DSL,37.245505,-118.06294299999999,1,98.9,0,8,None,1826,0,0,1,0,58,1,0.0,1804.38,0.0,5780.7,0,1,93513
4051,0,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),97.7,6869.7,0,26,58,28.59,5406,0,Bishop,0,0,Fiber Optic,37.045840000000005,-118.397236,1,97.7,0,7,Offer A,13309,0,0,1,1,72,1,3984.0,2058.48,0.0,6869.7,1,0,93514
4052,0,1,0,0,30,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,40.3,1172.95,1,74,8,0.0,3016,1,Boron,1,0,Cable,34.957029999999996,-117.73045,0,41.912,0,0,None,2241,0,0,0,0,30,0,0.0,0.0,0.0,1172.95,0,1,93516
4053,1,1,0,0,11,1,1,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),60.25,662.95,0,75,17,48.33,5296,0,Bridgeport,0,1,DSL,38.184583,-119.28655800000001,0,60.25,0,0,None,826,0,0,0,0,11,2,0.0,531.63,0.0,662.95,0,1,93517
4054,0,1,0,0,34,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,56.25,1765.95,0,72,28,0.0,5597,0,Caliente,1,0,Fiber Optic,35.358953,-118.527064,0,56.25,0,0,None,1022,0,1,0,0,34,1,494.0,0.0,0.0,1765.95,0,0,93518
4055,1,0,0,0,54,0,No phone service,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),46.2,2431.95,0,51,7,0.0,6143,0,Darwin,0,1,Cable,36.319181,-117.593053,0,46.2,0,0,Offer B,64,0,0,0,1,54,1,0.0,0.0,0.0,2431.95,0,1,93522
4056,0,0,0,0,3,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,50.6,155.35,1,56,28,0.0,4800,1,Edwards,0,0,Cable,34.966777,-117.961179,0,52.623999999999995,0,0,None,7685,0,0,0,1,3,1,0.0,0.0,0.0,155.35,0,1,93523
4057,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.9,1859.2,0,42,0,18.21,5192,0,Independence,0,0,NA,36.869584,-118.189241,1,24.9,3,5,Offer A,734,0,0,1,0,72,2,0.0,1311.12,0.0,1859.2,0,0,93526
4058,0,0,1,1,40,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,84.85,3303.05,1,64,21,2.03,5764,1,Temecula,1,0,DSL,33.507255,-117.029473,1,88.244,0,1,Offer B,46171,1,0,1,0,40,3,694.0,81.19999999999997,0.0,3303.05,0,0,92592
4059,0,0,1,1,2,1,0,DSL,0,0,1,1,Month-to-month,0,Mailed check,65.7,134.35,1,21,56,27.27,4265,1,Johannesburg,0,0,DSL,35.363339,-117.63764099999999,1,68.328,2,1,None,207,0,1,1,1,2,1,75.0,54.54,0.0,134.35,1,0,93528
4060,1,0,1,1,54,1,1,DSL,0,0,0,1,Two year,0,Credit card (automatic),63.35,3409.1,0,29,59,36.09,4232,0,June Lake,1,1,Fiber Optic,37.730269,-119.05581299999999,1,63.35,3,1,Offer B,618,0,0,1,1,54,0,0.0,1948.86,0.0,3409.1,1,1,93529
4061,0,0,0,0,14,1,0,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),50.1,709.5,0,19,59,36.22,2331,0,Keeler,0,0,Cable,36.560497999999995,-117.962461,0,50.1,0,0,None,71,0,0,0,0,14,1,419.0,507.08,0.0,709.5,1,0,93530
4062,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.5,70.5,1,53,3,41.39,4123,1,Keene,0,0,DSL,35.214982,-118.59048999999999,0,73.32000000000002,0,0,None,1436,0,0,0,0,1,3,0.0,41.39,0.0,70.5,0,0,93531
4063,0,0,0,0,10,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,94.85,953.45,1,34,23,43.26,3074,1,Lake Hughes,1,0,Cable,34.659579,-118.58421200000001,0,98.644,0,0,None,2771,0,0,0,1,10,4,219.0,432.6,0.0,953.45,0,0,93532
4064,0,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,50.15,50.15,0,63,24,38.33,4421,0,Lancaster,0,0,Fiber Optic,34.727529,-118.153098,0,50.15,0,0,Offer E,35109,0,0,0,0,1,0,0.0,38.33,0.0,50.15,0,1,93534
4065,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.75,19.75,1,21,0,29.33,4851,1,Lancaster,0,1,NA,34.712708,-117.889656,0,19.75,0,0,None,57794,0,1,0,0,1,2,0.0,29.33,0.0,19.75,1,0,93535
4066,1,0,0,0,56,1,1,DSL,1,1,0,0,One year,1,Bank transfer (automatic),64.65,3665.55,0,22,59,48.32,4656,0,Lancaster,0,1,Fiber Optic,34.741406,-118.38111,0,64.65,0,0,Offer B,49309,1,0,0,0,56,1,2163.0,2705.92,0.0,3665.55,1,0,93536
4067,0,0,1,0,68,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),79.6,5515.8,0,38,14,47.95,5601,0,Lee Vining,0,0,DSL,37.890145000000004,-119.184087,1,79.6,0,7,Offer A,504,1,0,1,1,68,0,0.0,3260.600000000001,0.0,5515.8,0,1,93541
4068,0,0,1,1,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.5,272,0,58,0,41.05,2993,0,Littlerock,0,0,NA,34.505272999999995,-117.955054,1,19.5,1,2,None,11198,0,0,1,0,14,2,0.0,574.6999999999998,0.0,272.0,0,0,93543
4069,1,0,1,1,68,1,0,Fiber optic,1,0,1,1,Two year,1,Electronic check,99.55,6668,0,38,28,38.75,4319,0,Llano,0,1,DSL,34.500091,-117.76586200000001,1,99.55,3,9,Offer A,1220,1,0,1,1,68,0,1867.0,2635.0,0.0,6668.0,0,0,93544
4070,1,1,1,0,55,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.0,4052.4,0,68,27,42.9,4958,0,Fallbrook,0,1,Fiber Optic,33.362575,-117.299644,1,74.0,0,6,None,42239,0,0,1,0,55,0,0.0,2359.5,0.0,4052.4,0,1,92028
4071,0,0,0,0,16,0,No phone service,DSL,1,0,1,0,Month-to-month,1,Electronic check,38.9,664.4,0,34,30,0.0,3300,0,Mammoth Lakes,0,0,DSL,37.550074,-118.837167,0,38.9,0,0,None,8217,0,0,0,0,16,0,199.0,0.0,0.0,664.4,0,0,93546
4072,1,1,0,0,9,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.55,718.55,0,73,15,24.85,5811,0,Olancha,0,1,Fiber Optic,36.296851000000004,-117.86546899999999,0,79.55,0,0,Offer E,318,0,0,0,0,9,3,0.0,223.65,0.0,718.55,0,1,93549
4073,1,0,1,1,14,1,0,DSL,1,1,1,0,Month-to-month,1,Electronic check,65.45,937.6,1,42,21,45.6,2881,1,Palmdale,0,1,Cable,34.536232,-118.082935,1,68.06800000000001,1,1,None,67232,0,3,1,0,14,3,0.0,638.4,0.0,937.6,0,1,93550
4074,1,1,1,0,58,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.7,5812.6,1,67,6,3.18,4662,1,Palmdale,1,1,Fiber Optic,34.613476,-118.256358,1,102.648,0,1,Offer B,34045,0,2,1,1,58,1,349.0,184.44,0.0,5812.6,0,0,93551
4075,1,0,0,0,53,0,No phone service,DSL,1,1,0,1,Month-to-month,1,Bank transfer (automatic),46.3,2546.85,0,37,24,0.0,6245,0,Palmdale,0,1,Fiber Optic,34.557711,-118.02944099999999,0,46.3,0,0,Offer B,25370,0,0,0,1,53,2,0.0,0.0,0.0,2546.85,0,1,93552
4076,1,0,1,0,70,1,1,Fiber optic,1,1,1,0,Two year,1,Credit card (automatic),99.35,6944.5,0,58,13,48.0,4120,0,Pearblossom,1,1,Fiber Optic,34.445239,-117.89486799999999,1,99.35,0,10,Offer A,1613,0,0,1,0,70,1,903.0,3360.0,0.0,6944.5,0,0,93553
4077,0,1,1,1,14,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.8,1346.3,0,79,30,14.39,3471,0,Randsburg,0,0,Cable,35.405722,-117.773354,1,95.8,1,5,None,117,0,0,1,0,14,1,404.0,201.46,0.0,1346.3,0,0,93554
4078,1,0,1,1,22,1,0,DSL,1,0,1,0,One year,1,Bank transfer (automatic),67.5,1544.05,1,49,19,19.8,3378,1,Temecula,1,1,DSL,33.507255,-117.029473,1,70.2,0,1,None,46171,1,0,1,0,22,5,0.0,435.6,0.0,1544.05,0,1,92592
4079,0,0,1,0,10,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),78.15,765.15,0,23,42,38.03,3403,0,Rosamond,0,0,Fiber Optic,34.903052,-118.41125100000001,1,78.15,0,4,None,14931,0,0,1,0,10,0,0.0,380.3,0.0,765.15,1,1,93560
4080,0,0,1,1,29,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,26.1,692.55,0,62,0,5.35,2828,0,Tehachapi,0,0,NA,35.073777,-118.65211200000002,1,26.1,2,8,None,25805,0,0,1,0,29,1,0.0,155.14999999999995,0.0,692.55,0,0,93561
4081,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.6,69.6,1,25,65,14.19,2412,1,Temecula,0,0,Cable,33.507255,-117.029473,0,72.384,0,0,None,46171,0,0,0,1,1,6,0.0,14.19,0.0,69.6,1,0,92592
4082,1,0,1,0,49,1,1,DSL,1,0,1,1,One year,0,Electronic check,84.35,4059.35,1,61,11,39.55,6452,1,Valyermo,1,1,Cable,34.39583,-117.734568,1,87.72399999999999,0,1,Offer B,413,1,2,1,1,49,3,447.0,1937.95,0.0,4059.35,0,0,93563
4083,0,1,1,0,68,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.2,6851.65,1,74,26,21.33,4481,1,Palmdale,0,0,Fiber Optic,34.598221,-117.79593,1,104.208,0,1,None,6787,0,0,1,1,68,1,1781.0,1450.4399999999996,0.0,6851.65,0,0,93591
4084,0,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,78.05,78.05,1,20,65,29.41,3458,1,Ahwahnee,0,0,Cable,37.375816,-119.739935,0,81.172,0,0,None,1968,0,0,0,1,1,3,0.0,29.41,0.0,78.05,1,1,93601
4085,0,0,0,0,30,0,No phone service,DSL,0,0,0,1,One year,1,Credit card (automatic),40.35,1187.05,0,23,42,0.0,5455,0,Auberry,0,0,Cable,36.991762,-119.242874,0,40.35,0,0,None,3464,1,0,0,1,30,1,0.0,0.0,0.0,1187.05,1,1,93602
4086,0,0,1,0,72,1,1,DSL,1,1,1,0,Two year,0,Credit card (automatic),79.2,5401.9,0,21,59,22.41,4288,0,Badger,1,0,DSL,36.64545,-118.924982,1,79.2,0,9,Offer A,273,1,0,1,0,72,2,0.0,1613.52,0.0,5401.9,1,1,93603
4087,0,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.9,247,0,27,0,12.39,4905,0,Bass Lake,0,0,NA,37.458366999999996,-119.34501100000001,0,20.9,0,0,None,613,0,0,0,0,10,2,0.0,123.9,0.0,247.0,1,0,93604
4088,1,0,0,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,73.6,520,1,63,31,38.07,2679,1,Big Creek,0,1,Cable,37.17277,-119.2997,0,76.544,0,0,None,273,0,0,0,0,7,2,161.0,266.49,0.0,520.0,0,0,93605
4089,0,0,0,0,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.75,706.6,1,55,13,16.48,5003,1,Biola,0,0,DSL,36.798882,-120.01951100000001,0,77.74000000000002,0,0,Offer E,807,0,2,0,0,9,2,92.0,148.32,0.0,706.6,0,0,93606
4090,0,0,0,1,1,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,49.9,49.9,0,39,53,9.0,5969,0,Cantua Creek,0,0,Fiber Optic,36.488056,-120.40769099999999,0,49.9,3,0,Offer E,1766,0,0,0,0,1,1,0.0,9.0,0.0,49.9,0,0,93608
4091,0,0,0,0,20,1,1,DSL,0,1,0,1,Month-to-month,1,Credit card (automatic),68.9,1370.35,0,44,11,22.75,3265,0,Caruthers,0,0,Fiber Optic,36.5276,-119.865999,0,68.9,0,0,None,5446,1,0,0,1,20,1,151.0,455.0,0.0,1370.35,0,0,93609
4092,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.25,20.25,0,42,0,28.18,5854,0,Chowchilla,0,0,NA,37.100947999999995,-120.27013600000001,0,20.25,0,0,Offer E,19391,0,0,0,0,1,1,0.0,28.18,0.0,20.25,0,0,93610
4093,0,0,0,0,29,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),76.0,2215.25,0,24,42,7.01,5324,0,Clovis,0,0,Cable,36.917652000000004,-119.59375700000001,0,76.0,0,0,None,46858,0,0,0,0,29,1,0.0,203.29,0.0,2215.25,1,1,93611
4094,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,74.0,74,0,34,25,23.7,4148,0,Clovis,0,1,DSL,36.814539,-119.711868,0,74.0,0,0,Offer E,33856,1,0,0,0,1,0,0.0,23.7,0.0,74.0,0,0,93612
4095,1,0,0,0,3,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,82.3,214.4,0,61,16,44.97,5755,0,Coarsegold,0,1,Fiber Optic,37.212191,-119.749323,0,82.3,0,0,None,9395,1,2,0,0,3,1,0.0,134.91,0.0,214.4,0,1,93614
4096,0,0,0,0,20,1,0,Fiber optic,1,0,1,0,Month-to-month,1,Bank transfer (automatic),89.4,1871.15,0,48,21,30.52,2098,0,Cutler,1,0,Fiber Optic,36.497895,-119.28548400000001,0,89.4,0,0,None,5519,0,0,0,0,20,0,393.0,610.4,0.0,1871.15,0,0,93615
4097,1,0,0,1,64,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),99.15,6171.2,0,31,24,22.41,4590,0,Del Rey,0,1,Cable,36.657462,-119.595293,0,99.15,1,0,Offer B,1965,1,0,0,1,64,0,1481.0,1434.24,0.0,6171.2,0,0,93616
4098,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.2,20.2,1,38,0,45.49,5355,1,Dinuba,0,1,NA,36.523619000000004,-119.38686799999999,0,20.2,0,0,Offer E,24206,0,0,0,0,1,2,0.0,45.49,0.0,20.2,0,0,93618
4099,0,0,0,0,6,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),29.45,161.45,0,22,52,0.0,4391,0,Dos Palos,0,0,DSL,37.045728000000004,-120.63068200000001,0,29.45,0,0,Offer E,9388,0,0,0,0,6,0,84.0,0.0,0.0,161.45,1,0,93620
4100,1,0,1,0,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,19.8,1013.2,0,55,0,1.87,5914,0,Dunlap,0,1,NA,36.789213000000004,-119.14033799999999,1,19.8,0,5,Offer B,506,0,0,1,0,50,1,0.0,93.5,0.0,1013.2,0,0,93621
4101,1,0,0,0,6,1,0,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),59.15,336.7,0,60,5,20.11,3613,0,Firebaugh,0,1,Fiber Optic,36.785618,-120.625382,0,59.15,0,0,Offer E,9491,0,0,0,1,6,0,1.68,120.66,0.0,336.7,0,1,93622
4102,1,0,1,1,7,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.75,333.65,0,42,17,28.7,4699,0,Fish Camp,0,1,Fiber Optic,37.483534999999996,-119.679414,1,44.75,1,7,Offer E,77,0,1,1,0,7,1,57.0,200.9,0.0,333.65,0,0,93623
4103,1,0,1,1,72,1,1,Fiber optic,0,0,0,1,Two year,1,Credit card (automatic),90.8,6511.8,0,22,59,23.7,6188,0,Five Points,1,1,DSL,36.397745,-120.11991100000002,1,90.8,1,1,Offer A,1852,0,0,1,1,72,0,384.2,1706.4,0.0,6511.8,1,1,93624
4104,1,0,1,0,8,1,0,DSL,0,1,0,0,Month-to-month,1,Bank transfer (automatic),49.55,393.45,0,24,53,2.38,5922,0,Fowler,0,1,Cable,36.625792,-119.67248300000001,1,49.55,0,6,Offer E,5635,0,0,1,0,8,1,209.0,19.04,0.0,393.45,1,0,93625
4105,0,0,1,1,67,1,1,Fiber optic,1,0,1,1,Two year,0,Credit card (automatic),106.7,7009.5,0,35,16,40.35,4780,0,Friant,0,0,DSL,37.027663000000004,-119.69056,1,106.7,2,3,Offer A,1125,1,0,1,1,67,1,0.0,2703.4500000000007,0.0,7009.5,0,1,93626
4106,0,1,1,0,24,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.55,2264.05,1,69,13,13.38,4937,1,Helm,0,0,DSL,36.520537,-120.118055,1,97.292,0,1,None,152,0,0,1,1,24,3,294.0,321.12,0.0,2264.05,0,0,93627
4107,0,0,1,0,72,1,1,Fiber optic,1,1,0,1,Two year,1,Credit card (automatic),94.45,6921.7,0,22,48,22.74,5274,0,Hume,0,0,Cable,36.807595,-118.901544,1,94.45,0,5,Offer A,93,0,0,1,1,72,0,3322.0,1637.28,0.0,6921.7,1,0,93628
4108,1,0,1,1,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.45,600.25,0,25,0,5.86,3470,0,Kerman,0,1,NA,36.727418,-120.123526,1,19.45,1,6,None,14062,0,0,1,0,33,2,0.0,193.38,0.0,600.25,1,0,93630
4109,1,0,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,25.05,56.35,1,22,80,0.0,4810,1,Kingsburg,0,1,Cable,36.478239,-119.52136999999999,0,26.052000000000003,0,0,Offer E,14088,0,0,0,1,2,0,45.0,0.0,0.0,56.35,1,0,93631
4110,1,0,1,0,70,1,0,DSL,1,1,0,1,Two year,0,Mailed check,67.95,4664.15,0,41,15,24.93,5514,0,Lakeshore,0,1,Fiber Optic,37.290606,-119.216328,1,67.95,0,7,Offer A,52,1,0,1,1,70,2,0.0,1745.1,0.0,4664.15,0,1,93634
4111,0,0,0,0,22,1,0,DSL,0,1,1,0,One year,0,Bank transfer (automatic),65.25,1441.8,0,22,85,1.74,5146,0,Los Banos,1,0,Fiber Optic,36.995162,-120.955099,0,65.25,0,0,None,29124,0,0,0,0,22,0,0.0,38.28,0.0,1441.8,1,1,93635
4112,0,0,0,0,59,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Bank transfer (automatic),99.45,5623.7,0,54,12,39.42,5247,0,Madera,1,0,Cable,36.902954,-120.194274,0,99.45,0,0,Offer B,28434,0,0,0,1,59,0,0.0,2325.78,0.0,5623.7,0,1,93637
4113,1,0,0,0,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.35,695.85,0,37,0,12.72,3526,0,Madera,0,1,NA,37.004068,-119.930027,0,20.35,0,0,None,49247,0,2,0,0,36,1,0.0,457.92,0.0,695.85,0,0,93638
4114,0,0,1,1,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.95,1028.75,0,60,0,14.54,4057,0,Escondido,0,0,NA,33.141265000000004,-116.967221,1,19.95,1,10,Offer B,48690,0,0,1,0,51,2,0.0,741.54,0.0,1028.75,0,0,92027
4115,1,0,1,0,53,1,1,DSL,1,0,1,0,One year,0,Bank transfer (automatic),77.4,4155.95,0,52,13,47.55,5313,0,Miramonte,1,1,Cable,36.696759,-119.024051,1,77.4,0,1,Offer B,571,1,0,1,0,53,0,0.0,2520.15,0.0,4155.95,0,1,93641
4116,0,0,1,1,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.7,395.6,0,50,0,7.31,4910,0,North Fork,0,0,NA,37.244307,-119.470256,1,19.7,3,7,None,3376,0,0,1,0,20,1,0.0,146.2,0.0,395.6,0,0,93643
4117,1,0,1,0,63,1,0,Fiber optic,1,0,1,1,Two year,0,Credit card (automatic),99.7,6330.4,0,46,6,26.81,5135,0,Oakhurst,1,1,DSL,37.648647,-119.231447,1,99.7,0,3,Offer B,8521,0,0,1,1,63,0,0.0,1689.03,0.0,6330.4,0,1,93644
4118,0,0,0,0,40,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Credit card (automatic),74.8,2971.7,0,50,15,18.57,3258,0,O Neals,0,0,Cable,37.140104,-119.65709199999999,0,74.8,0,0,Offer B,173,0,0,0,0,40,1,0.0,742.8,0.0,2971.7,0,1,93645
4119,1,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.15,638,0,53,0,7.74,4052,0,Orange Cove,0,1,NA,36.633497999999996,-119.298895,0,19.15,0,0,None,8449,0,0,0,0,35,1,0.0,270.90000000000003,0.0,638.0,0,0,93646
4120,1,0,1,1,26,1,0,Fiber optic,0,0,0,1,One year,0,Bank transfer (automatic),78.95,2034.25,0,54,75,24.17,4237,0,Orosi,0,1,Cable,36.600184999999996,-119.175655,1,78.95,3,3,None,9780,0,0,1,1,26,0,0.0,628.4200000000002,0.0,2034.25,0,1,93647
4121,1,1,1,0,27,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,95.55,2510.2,1,70,8,39.49,2999,1,Parlier,1,1,DSL,36.622237,-119.521126,1,99.37200000000001,0,1,None,12587,0,1,1,1,27,2,201.0,1066.23,0.0,2510.2,0,0,93648
4122,1,0,0,1,53,1,0,DSL,1,1,0,0,One year,0,Credit card (automatic),62.85,3419.5,0,20,59,47.81,6281,0,Fresno,0,1,Fiber Optic,36.841654999999996,-119.79711299999998,0,62.85,2,0,Offer B,3258,1,0,0,0,53,0,2018.0,2533.9300000000007,0.0,3419.5,1,0,93650
4123,1,1,1,0,34,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),71.55,2427.35,0,72,8,12.98,3583,0,Prather,0,1,DSL,37.007238,-119.505661,1,71.55,0,2,None,1314,0,1,1,0,34,2,194.0,441.32,0.0,2427.35,0,0,93651
4124,0,1,1,0,19,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.95,1760.25,0,78,27,19.57,5316,0,Raisin City,0,0,Cable,36.594542,-119.905245,1,94.95,0,10,None,265,0,0,1,0,19,2,0.0,371.83,0.0,1760.25,0,1,93652
4125,1,0,1,0,43,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),86.1,3551.65,0,48,20,7.63,2358,0,Raymond,1,1,Fiber Optic,37.252057,-119.95783,1,86.1,0,10,Offer B,972,0,0,1,0,43,1,71.03,328.09,0.0,3551.65,0,1,93653
4126,1,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.55,122.9,0,48,0,36.54,3072,0,Reedley,0,1,NA,36.636638,-119.421842,1,19.55,3,5,Offer E,25923,0,0,1,0,6,0,0.0,219.24,0.0,122.9,0,0,93654
4127,1,0,0,1,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.8,1424.2,0,48,0,22.47,4262,0,Riverdale,0,1,NA,36.452211,-119.94575,0,24.8,3,0,Offer B,5729,0,1,0,0,56,1,0.0,1258.32,0.0,1424.2,0,0,93656
4128,1,0,0,0,57,0,No phone service,DSL,0,1,1,0,Month-to-month,1,Electronic check,39.3,2111.45,1,23,65,0.0,4917,1,Sanger,0,1,DSL,36.819628,-119.44041399999999,0,40.872,0,0,Offer B,28991,0,0,0,1,57,6,1372.0,0.0,0.0,2111.45,1,0,93657
4129,1,0,1,1,34,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,84.05,2909.95,0,63,26,5.65,3476,0,San Joaquin,1,1,Fiber Optic,36.600193,-120.153393,1,84.05,1,10,None,4318,0,0,1,0,34,2,0.0,192.1,0.0,2909.95,0,1,93660
4130,0,0,0,0,10,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,36.25,374,0,33,23,0.0,4571,0,Selma,0,0,Fiber Optic,36.545322,-119.64228100000001,0,36.25,0,0,None,26213,1,0,0,0,10,0,86.0,0.0,0.0,374.0,0,0,93662
4131,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.25,20.25,1,64,0,10.71,2783,1,Shaver Lake,0,0,NA,37.223,-119.001021,0,20.25,0,0,Offer E,642,0,0,0,0,1,2,0.0,10.71,0.0,20.25,0,0,93664
4132,0,0,0,0,13,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,23.9,300.8,1,30,58,0.0,2967,1,South Dos Palos,0,0,DSL,36.959731,-120.65351899999999,0,24.856,0,0,None,343,0,0,0,0,13,3,174.0,0.0,0.0,300.8,0,0,93665
4133,1,0,0,0,56,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,98.6,5581.05,0,62,28,10.99,5601,0,Sultana,0,1,Fiber Optic,36.545353000000006,-119.33853500000001,0,98.6,0,0,Offer B,306,0,0,0,1,56,1,0.0,615.44,0.0,5581.05,0,1,93666
4134,0,0,1,0,55,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),103.65,5676.65,0,54,25,33.66,4768,0,Tollhouse,1,0,Cable,36.993666,-119.34826699999999,1,103.65,0,4,Offer B,2633,0,0,1,1,55,2,0.0,1851.3,0.0,5676.65,0,1,93667
4135,0,0,1,1,36,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),92.9,3379.25,0,23,59,40.54,3570,0,Tranquillity,1,0,Fiber Optic,36.635661,-120.28864399999999,1,92.9,2,7,None,1130,1,0,1,1,36,1,0.0,1459.44,0.0,3379.25,1,1,93668
4136,1,0,1,0,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.9,942.95,0,26,0,43.2,5394,0,Wishon,0,1,NA,37.287758000000004,-119.548156,1,19.9,0,0,Offer B,327,0,0,0,0,47,0,0.0,2030.4,0.0,942.95,1,0,93669
4137,0,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.1,232.4,0,43,0,24.65,2360,0,Traver,0,0,NA,36.456091,-119.486225,1,20.1,1,3,None,646,0,0,1,0,12,0,0.0,295.7999999999999,0.0,232.4,0,0,93673
4138,0,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.45,85.45,1,48,25,22.97,4931,1,Squaw Valley,1,0,Cable,36.719141,-119.20267700000001,0,88.86800000000002,0,0,Offer E,3146,0,0,0,0,1,4,0.0,22.97,0.0,85.45,0,0,93675
4139,1,1,0,0,24,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.5,2088.45,0,76,23,46.13,4422,0,Fresno,0,1,Cable,36.749403,-119.78757399999999,0,80.5,0,0,None,13858,0,0,0,0,24,1,0.0,1107.12,0.0,2088.45,0,1,93701
4140,0,0,0,0,63,1,1,Fiber optic,0,1,1,1,One year,0,Bank transfer (automatic),99.9,6137,1,22,65,8.38,4776,1,Fresno,0,0,Cable,36.739385,-119.753649,0,103.89600000000002,0,0,Offer B,47999,0,0,0,1,63,1,3989.0,527.94,0.0,6137.0,1,0,93702
4141,0,1,0,0,35,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,39.85,1434.6,0,77,26,0.0,2030,0,Fresno,1,0,DSL,36.768774,-119.76263300000001,0,39.85,0,0,None,31180,0,1,0,0,35,1,373.0,0.0,0.0,1434.6,0,0,93703
4142,0,0,0,0,67,1,0,DSL,1,1,0,0,One year,0,Credit card (automatic),60.5,3870,0,28,73,35.99,4363,0,Fresno,0,0,DSL,36.799648,-119.801247,0,60.5,0,0,Offer A,26580,1,0,0,0,67,0,282.51,2411.33,0.0,3870.0,1,1,93704
4143,1,0,0,0,25,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.8,2043.45,1,64,24,8.31,4203,1,Fresno,0,1,DSL,36.787240000000004,-119.82781299999999,0,88.19200000000001,0,0,Offer C,35451,0,1,0,1,25,1,490.0,207.75,0.0,2043.45,0,0,93705
4144,1,0,0,0,21,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Mailed check,103.85,2215,0,60,3,15.89,4520,0,Fresno,1,1,Fiber Optic,36.654614,-119.903674,0,103.85,0,0,Offer D,35790,0,0,0,1,21,3,0.0,333.69,0.0,2215.0,0,1,93706
4145,0,0,0,0,13,1,0,DSL,1,1,0,1,Month-to-month,0,Bank transfer (automatic),67.8,842.25,0,36,30,28.45,4115,0,Fresno,0,0,Cable,36.822715,-119.761826,0,67.8,0,0,Offer D,29337,1,0,0,1,13,0,0.0,369.85,0.0,842.25,0,1,93710
4146,1,0,1,0,35,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.2,2576.2,1,48,13,48.47,4639,1,San Dimas,0,1,Cable,34.102119,-117.815532,1,78.20800000000001,0,1,Offer C,33878,0,0,1,0,35,4,335.0,1696.45,0.0,2576.2,0,0,91773
4147,1,1,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.85,1901,0,69,0,22.19,4367,0,Fresno,0,1,NA,36.878709,-119.7645,1,24.85,0,0,Offer A,45087,0,0,0,0,71,0,0.0,1575.49,0.0,1901.0,0,0,93720
4148,0,0,0,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.35,601.6,0,46,0,2.76,5227,0,Fresno,0,0,NA,36.732694,-119.783786,0,19.35,0,0,None,6848,0,0,0,0,29,1,0.0,80.03999999999998,0.0,601.6,0,0,93721
4149,1,0,1,0,71,0,No phone service,DSL,0,1,1,1,Two year,0,Electronic check,49.35,3515.25,1,44,28,0.0,4879,1,Fresno,0,1,DSL,36.78979,-119.92989399999999,1,51.32400000000001,0,1,None,60889,0,1,1,1,71,1,984.0,0.0,0.0,3515.25,0,0,93722
4150,1,1,1,0,7,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.0,605.45,0,71,11,41.97,5711,0,Fresno,0,1,Cable,36.623632,-119.741322,1,89.0,0,8,None,21010,0,0,1,1,7,1,0.0,293.79,0.0,605.45,0,1,93725
4151,0,1,0,0,57,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,55.0,3094.05,0,65,26,0.0,4622,0,Fresno,1,0,Fiber Optic,36.793601,-119.761131,0,55.0,0,0,Offer B,39148,0,0,0,1,57,0,0.0,0.0,0.0,3094.05,0,1,93726
4152,1,0,1,0,65,1,1,DSL,1,0,0,1,Two year,0,Bank transfer (automatic),76.15,4929.55,0,45,13,21.58,6177,0,Fresno,1,1,Fiber Optic,36.751489,-119.68072,1,76.15,0,2,Offer B,54701,1,0,1,1,65,0,0.0,1402.6999999999996,0.0,4929.55,0,1,93727
4153,1,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.3,595.05,0,44,0,21.66,3159,0,Fresno,0,1,NA,36.757345,-119.818274,0,20.3,0,0,None,16346,0,0,0,0,27,0,0.0,584.82,0.0,595.05,0,0,93728
4154,1,0,0,0,6,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.9,469.8,1,49,12,6.32,4160,1,Salinas,0,1,DSL,36.64152,-121.622188,0,77.89600000000002,0,0,None,35739,0,3,0,0,6,2,56.0,37.92,0.0,469.8,0,0,93901
4155,0,1,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),117.35,8436.25,0,78,30,14.94,4008,0,Salinas,1,0,Cable,36.667794,-121.60130600000001,0,117.35,0,0,Offer A,58548,1,0,0,1,72,1,2531.0,1075.68,0.0,8436.25,0,0,93905
4156,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.75,19.75,0,31,0,10.22,4441,0,Salinas,0,1,NA,36.722898,-121.633648,0,19.75,0,0,Offer E,53946,0,0,0,0,1,1,0.0,10.22,0.0,19.75,0,0,93906
4157,1,0,0,0,11,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),45.2,492,0,44,22,40.59,5253,0,Salinas,0,1,DSL,36.77462,-121.66471399999999,0,45.2,0,0,Offer D,22292,0,0,0,0,11,0,108.0,446.49,0.0,492.0,0,0,93907
4158,1,0,1,1,39,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.2,987.95,0,64,0,20.49,5453,0,Salinas,0,1,NA,36.624338,-121.615669,1,25.2,2,8,None,13027,0,0,1,0,39,1,0.0,799.1099999999999,0.0,987.95,0,0,93908
4159,0,1,0,0,59,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,89.75,5496.9,0,80,5,25.57,5170,0,Escondido,1,0,Fiber Optic,33.141265000000004,-116.967221,0,89.75,0,0,Offer B,48690,0,0,0,0,59,0,275.0,1508.63,0.0,5496.9,0,0,92027
4160,1,0,0,0,26,1,0,DSL,1,0,1,1,One year,0,Bank transfer (automatic),75.0,1908.35,0,24,76,49.61,4705,0,Carmel By The Sea,0,1,DSL,36.554618,-121.92223899999999,0,75.0,0,0,None,2966,1,0,0,1,26,2,0.0,1289.86,0.0,1908.35,1,1,93921
4161,1,1,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,49.95,107.1,0,71,9,37.97,5251,0,Carmel,1,1,DSL,36.460611,-121.852507,0,49.95,0,0,Offer E,13121,0,0,0,0,2,1,0.0,75.94,0.0,107.1,0,1,93923
4162,0,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),65.7,4575.35,0,44,23,0.0,6187,0,Carmel Valley,1,0,DSL,36.414611,-121.6386,1,65.7,2,5,Offer A,6691,1,0,1,1,72,0,1052.0,0.0,0.0,4575.35,0,0,93924
4163,1,0,1,0,65,1,1,DSL,1,1,0,0,One year,0,Credit card (automatic),67.05,4309.55,0,50,18,39.49,5224,0,Chualar,1,1,Fiber Optic,36.596271,-121.442274,1,67.05,0,6,Offer B,1140,0,0,1,0,65,0,776.0,2566.85,0.0,4309.55,0,0,93925
4164,1,0,1,1,72,1,1,Fiber optic,0,1,1,1,Two year,0,Credit card (automatic),110.9,7922.75,0,31,11,45.32,6444,0,Gonzales,1,1,Fiber Optic,36.52588,-121.39671899999999,1,110.9,1,5,Offer A,9023,1,0,1,1,72,1,872.0,3263.04,0.0,7922.75,0,0,93926
4165,1,0,0,0,6,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),87.95,522.35,0,37,12,43.37,2684,0,Greenfield,0,1,Fiber Optic,36.248708,-121.38661699999999,0,87.95,0,0,None,14204,1,0,0,1,6,0,63.0,260.22,0.0,522.35,0,0,93927
4166,1,1,0,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.8,587.7,0,79,0,25.89,3836,0,Jolon,0,1,NA,35.930782,-121.189757,0,19.8,0,0,None,254,0,0,0,0,32,0,0.0,828.48,0.0,587.7,0,0,93928
4167,0,0,1,0,50,1,1,DSL,0,0,1,1,One year,0,Bank transfer (automatic),75.7,3876.2,0,40,28,9.47,6144,0,King City,1,0,Fiber Optic,36.220760999999996,-120.980777,1,75.7,0,5,Offer B,14477,0,1,1,1,50,2,1085.0,473.50000000000006,0.0,3876.2,0,0,93930
4168,1,0,1,0,61,0,No phone service,DSL,1,0,1,1,Two year,1,Mailed check,62.15,3778.85,0,22,59,0.0,6427,0,Lockwood,1,1,Fiber Optic,35.989792,-121.05593300000001,1,62.15,0,1,Offer B,538,1,0,1,1,61,0,0.0,0.0,0.0,3778.85,1,1,93932
4169,0,0,0,0,15,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.25,1457.25,1,43,29,16.82,3968,1,Marina,1,0,Fiber Optic,36.689582,-121.758398,0,105.3,0,0,None,21759,0,0,0,1,15,3,423.0,252.3,0.0,1457.25,0,0,93933
4170,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),115.15,8349.45,0,29,58,35.71,5398,0,Monterey,1,1,DSL,36.362741,-121.869685,1,115.15,0,4,Offer A,32857,1,0,1,1,72,3,0.0,2571.12,0.0,8349.45,1,1,93940
4171,1,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,18.95,185.6,1,59,0,49.74,5403,1,Pacific Grove,0,1,NA,36.618337,-121.92641699999999,0,18.95,0,0,Offer E,15449,0,1,0,0,9,2,0.0,447.66,0.0,185.6,0,0,93950
4172,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.5,19.5,0,42,0,20.11,3107,0,Pebble Beach,0,0,NA,36.587497,-121.94481499999999,0,19.5,0,0,Offer E,4602,0,0,0,0,1,0,0.0,20.11,0.0,19.5,0,0,93953
4173,0,0,0,0,12,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.55,1066.9,0,33,25,18.75,2061,0,San Lucas,0,0,DSL,36.125529,-120.864443,0,86.55,0,0,Offer D,521,0,0,0,1,12,2,267.0,225.0,0.0,1066.9,0,0,93954
4174,0,0,0,0,37,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),28.6,973.55,1,31,11,0.0,4429,1,Seaside,0,0,DSL,36.625114,-121.82356499999999,0,29.744000000000003,0,0,None,38244,1,0,0,0,37,2,107.0,0.0,0.0,973.55,0,0,93955
4175,1,0,1,1,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.4,1226.45,0,42,0,31.49,5897,0,Soledad,0,1,NA,36.414215999999996,-121.360597,1,20.4,3,7,Offer B,13003,0,1,1,0,61,1,0.0,1920.89,0.0,1226.45,0,0,93960
4176,1,0,1,1,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.8,342.3,0,39,0,45.18,4808,0,Spreckels,0,1,NA,36.624641,-121.647195,1,19.8,3,1,Offer D,407,0,0,1,0,18,0,0.0,813.24,0.0,342.3,0,0,93962
4177,1,0,0,1,21,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.65,985.05,0,60,29,19.57,5731,0,Belmont,0,1,Fiber Optic,37.509366,-122.306132,0,45.65,2,0,Offer D,25566,0,0,0,0,21,1,0.0,410.97,0.0,985.05,0,1,94002
4178,1,0,1,1,68,0,No phone service,DSL,1,1,0,1,Two year,1,Mailed check,56.4,3948.45,0,47,19,0.0,4556,0,Brisbane,1,1,DSL,37.684694,-122.40711999999999,1,56.4,2,10,Offer A,3635,1,0,1,1,68,1,750.0,0.0,0.0,3948.45,0,0,94005
4179,1,1,0,0,12,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),73.3,828.05,0,78,24,43.4,5159,0,Burlingame,0,1,Fiber Optic,37.57028,-122.365778,0,73.3,0,0,None,40346,0,0,0,0,12,1,0.0,520.8,0.0,828.05,0,1,94010
4180,0,1,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,24.35,41.85,1,79,12,0.0,3278,1,Daly City,0,0,DSL,37.691561,-122.445202,0,25.324,0,0,None,47453,0,0,0,0,2,0,5.0,0.0,0.0,41.85,0,0,94014
4181,0,0,1,0,62,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.35,6164.7,0,30,82,15.06,5049,0,Daly City,1,0,Fiber Optic,37.680844,-122.48131000000001,1,101.35,0,10,Offer B,63337,0,0,1,1,62,0,0.0,933.72,0.0,6164.7,0,1,94015
4182,0,1,0,0,29,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,98.65,2862.75,1,76,18,20.98,4235,1,Half Moon Bay,0,0,Cable,37.45567,-122.407992,0,102.596,0,0,None,17929,1,0,0,0,29,3,515.0,608.42,0.0,2862.75,0,0,94019
4183,1,0,0,1,1,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Mailed check,33.6,33.6,0,44,19,0.0,4369,0,La Honda,0,1,Fiber Optic,37.285677,-122.22416499999999,0,33.6,1,0,Offer E,1622,1,0,0,0,1,2,0.0,0.0,0.0,33.6,0,0,94020
4184,1,1,1,0,5,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),79.9,343.95,1,78,15,6.66,4324,1,Loma Mar,1,1,Fiber Optic,37.266388,-122.26308,1,83.096,0,1,None,148,0,0,1,0,5,2,52.0,33.3,0.0,343.95,0,0,94021
4185,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.7,20.7,0,27,0,45.86,3061,0,Los Altos,0,0,NA,37.349546000000004,-122.13435600000001,0,20.7,0,0,None,18486,0,0,0,0,1,0,0.0,45.86,0.0,20.7,1,0,94022
4186,1,0,0,1,62,1,1,Fiber optic,0,0,1,1,Two year,1,Electronic check,104.05,6590.5,0,44,19,17.67,5900,0,Los Altos,1,1,Cable,37.352911,-122.093002,0,104.05,1,0,Offer B,21496,1,1,0,1,62,1,0.0,1095.5400000000004,0.0,6590.5,0,1,94024
4187,0,0,1,1,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.25,717.95,0,26,0,42.51,5272,0,Menlo Park,0,0,NA,37.449551,-122.18376200000002,1,20.25,2,8,Offer C,39062,0,0,1,0,36,0,0.0,1530.36,0.0,717.95,1,0,94025
4188,0,1,0,0,28,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,103.3,2890.65,1,79,11,28.14,4136,1,Atherton,1,0,Fiber Optic,37.454924,-122.20316799999999,0,107.432,0,0,None,6876,1,1,0,0,28,5,318.0,787.9200000000002,0.0,2890.65,0,0,94027
4189,0,0,1,1,69,1,1,DSL,1,1,1,0,One year,0,Credit card (automatic),73.7,4885.85,0,59,21,7.84,4268,0,Portola Valley,0,0,Fiber Optic,37.369709,-122.21584399999999,1,73.7,3,10,Offer A,6601,1,0,1,0,69,1,1026.0,540.96,0.0,4885.85,0,0,94028
4190,0,0,1,0,11,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Credit card (automatic),96.2,1222.05,1,60,21,26.88,3101,1,Millbrae,0,0,Cable,37.601248,-122.403099,1,100.04799999999999,0,5,None,20350,1,2,1,0,11,3,0.0,295.68,0.0,1222.05,0,1,94030
4191,0,0,1,0,63,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,108.75,6871.7,0,49,26,20.37,4582,0,Montara,1,0,Fiber Optic,37.540582,-122.50959399999999,1,108.75,0,10,Offer B,2346,1,0,1,1,63,1,0.0,1283.3100000000004,0.0,6871.7,0,1,94037
4192,1,0,0,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.15,405.6,0,63,0,26.37,4402,0,Moss Beach,0,1,NA,37.515556,-122.502311,0,20.15,0,0,Offer D,3064,0,0,0,0,23,2,0.0,606.51,0.0,405.6,0,0,94038
4193,1,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.75,208.25,0,24,0,20.29,3926,0,Mountain View,0,1,NA,37.380662,-122.086022,0,19.75,0,0,Offer D,32143,0,1,0,0,10,2,0.0,202.9,0.0,208.25,1,0,94040
4194,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.95,1801.9,0,42,0,24.71,5072,0,Mountain View,0,0,NA,37.388349,-122.075299,1,25.95,0,2,Offer A,13483,0,0,1,0,71,0,0.0,1754.41,0.0,1801.9,0,0,94041
4195,0,1,0,0,45,1,1,DSL,1,0,0,1,Month-to-month,1,Electronic check,70.05,3062.45,0,80,3,18.46,4223,0,Mountain View,0,0,DSL,37.419725,-122.062947,0,70.05,0,0,Offer B,27822,1,0,0,1,45,0,92.0,830.7,0.0,3062.45,0,0,94043
4196,0,0,1,1,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.05,1764.75,0,24,0,4.27,4722,0,Pacifica,0,0,NA,37.573633,-122.45516699999999,1,24.05,2,4,Offer A,38885,0,0,1,0,70,0,0.0,298.9,0.0,1764.75,1,0,94044
4197,0,0,0,1,22,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.75,1816.75,0,32,19,33.73,4240,0,Pescadero,0,0,DSL,37.22565,-122.297533,0,84.75,2,0,Offer D,2055,0,0,0,1,22,0,345.0,742.06,0.0,1816.75,0,0,94060
4198,0,0,1,1,52,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,23.05,1255.1,0,42,0,19.21,4922,0,Redwood City,0,0,NA,37.461251000000004,-122.23541399999999,1,23.05,2,1,None,35737,0,0,1,0,52,1,0.0,998.92,0.0,1255.1,0,0,94061
4199,1,0,1,0,55,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,104.15,5743.05,1,21,84,10.61,4369,1,Redwood City,1,1,Fiber Optic,37.410567,-122.297152,1,108.31600000000002,0,1,Offer B,25569,1,2,1,1,55,4,4824.0,583.55,0.0,5743.05,1,0,94062
4200,0,0,0,0,65,0,No phone service,DSL,1,0,1,1,Two year,0,Credit card (automatic),59.95,3921.1,0,45,22,0.0,6251,0,Redwood City,1,0,Fiber Optic,37.499411,-122.19631799999999,0,59.95,0,0,None,32368,1,0,0,1,65,2,0.0,0.0,0.0,3921.1,0,1,94063
4201,0,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.55,1463.45,0,58,0,17.33,4424,0,Redwood City,0,0,NA,37.527497,-122.23094099999999,1,19.55,1,6,None,10658,0,0,1,0,72,1,0.0,1247.7599999999998,0.0,1463.45,0,0,94065
4202,1,0,1,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.6,189.45,0,23,0,39.35,3778,0,San Bruno,0,1,NA,37.624435999999996,-122.43066100000001,1,19.6,0,3,Offer D,39566,0,0,1,0,10,2,0.0,393.5,0.0,189.45,1,0,94066
4203,0,0,0,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.05,96.8,0,56,0,49.66,3810,0,San Carlos,0,0,NA,37.497915,-122.26736100000001,0,20.05,3,0,Offer E,28098,0,0,0,0,7,0,0.0,347.62,0.0,96.8,0,0,94070
4204,1,1,0,0,5,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,85.55,408.5,0,67,15,18.38,2850,0,San Gregorio,0,1,Cable,37.331762,-122.341444,0,85.55,0,0,Offer E,291,0,0,0,1,5,0,0.0,91.9,0.0,408.5,0,1,94074
4205,0,0,1,1,24,1,1,DSL,1,0,1,1,Two year,0,Credit card (automatic),78.6,1846.65,0,63,56,21.43,2939,0,South San Francisco,1,0,Cable,37.654436,-122.426468,1,78.6,3,8,Offer C,60599,0,0,1,1,24,0,0.0,514.3199999999998,0.0,1846.65,0,1,94080
4206,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),116.8,8456.75,0,25,59,16.01,6252,0,Sunnyvale,1,0,DSL,37.378541,-122.02045600000001,1,116.8,2,2,None,64010,1,0,1,1,72,0,498.95,1152.72,0.0,8456.75,1,1,94086
4207,1,0,0,0,21,0,No phone service,DSL,1,0,1,0,Month-to-month,1,Mailed check,43.55,1011.5,0,29,26,0.0,5808,0,Sunnyvale,0,1,DSL,37.3511,-122.03731100000002,0,43.55,0,0,Offer D,50070,1,2,0,0,21,1,0.0,0.0,0.0,1011.5,1,1,94087
4208,1,0,1,0,69,0,No phone service,DSL,0,1,1,1,One year,1,Credit card (automatic),60.8,4263.4,0,23,42,0.0,5683,0,Sunnyvale,1,1,Fiber Optic,37.421633,-122.00961299999999,1,60.8,0,7,None,16985,1,1,1,1,69,1,1791.0,0.0,0.0,4263.4,1,0,94089
4209,1,0,1,1,44,1,0,DSL,0,1,0,0,Month-to-month,1,Bank transfer (automatic),54.9,2549.1,0,58,52,46.54,4412,0,San Francisco,0,1,Cable,37.7795,-122.419233,1,54.9,3,4,None,28998,1,0,1,0,44,2,0.0,2047.76,0.0,2549.1,0,1,94102
4210,0,1,1,1,61,1,1,DSL,0,0,1,0,One year,1,Electronic check,65.2,3965.05,0,74,10,39.31,6238,0,San Francisco,1,0,DSL,37.773146999999994,-122.41128700000002,1,65.2,1,9,Offer B,23036,0,1,1,0,61,1,0.0,2397.9100000000008,0.0,3965.05,0,1,94103
4211,1,1,0,0,24,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),102.95,2496.7,1,73,29,3.23,5245,1,San Francisco,1,1,DSL,37.791222,-122.40224099999999,0,107.068,0,0,None,384,0,0,0,0,24,4,724.0,77.52,0.0,2496.7,0,0,94104
4212,0,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,90.6,90.6,1,41,24,31.68,2540,1,San Francisco,0,0,Fiber Optic,37.789168,-122.395009,0,94.22399999999999,0,0,Offer E,2066,0,0,0,1,1,4,0.0,31.68,0.0,90.6,0,0,94105
4213,0,0,0,0,6,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),50.8,288.05,1,51,13,21.91,4713,1,San Francisco,0,0,DSL,37.768881,-122.395521,0,52.832,0,0,Offer E,17372,1,1,0,0,6,2,3.74,131.46,0.0,288.05,0,1,94107
4214,1,0,0,0,4,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,90.05,368.1,1,42,12,12.24,3212,1,San Francisco,0,1,DSL,37.791998,-122.408653,0,93.652,0,0,Offer E,13723,0,0,0,1,4,1,44.0,48.96,0.0,368.1,0,0,94108
4215,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,108.2,7840.6,0,21,71,14.19,4773,0,San Francisco,1,1,DSL,37.794487,-122.42227,1,108.2,0,10,None,56330,1,0,1,1,72,2,0.0,1021.68,0.0,7840.6,1,1,94109
4216,1,0,0,0,72,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),92.0,6632.75,0,55,20,45.41,4200,0,San Francisco,1,1,DSL,37.750021000000004,-122.415201,0,92.0,0,0,None,74641,1,0,0,1,72,1,1327.0,3269.5199999999995,0.0,6632.75,0,0,94110
4217,1,1,1,0,14,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.1,1013.35,0,73,4,45.46,3771,0,San Francisco,0,1,DSL,37.801776000000004,-122.402293,1,75.1,0,8,None,3337,0,0,1,0,14,0,41.0,636.44,0.0,1013.35,0,0,94111
4218,1,0,0,0,7,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),25.05,152.95,0,26,0,45.13,4868,0,San Francisco,0,1,NA,37.720498,-122.443119,0,25.05,0,0,Offer E,73117,0,0,0,0,7,0,0.0,315.91,0.0,152.95,1,0,94112
4219,0,0,0,0,48,1,0,Fiber optic,0,1,0,0,One year,0,Electronic check,75.15,3772.65,0,64,23,41.26,3345,0,San Francisco,0,0,Fiber Optic,37.758084999999994,-122.43480100000001,0,75.15,0,0,None,30587,0,1,0,0,48,1,868.0,1980.48,0.0,3772.65,0,0,94114
4220,1,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.5,1026.35,0,43,0,36.23,5067,0,San Francisco,0,1,NA,37.786031,-122.437301,1,19.5,3,5,None,33122,0,0,1,0,55,3,0.0,1992.65,0.0,1026.35,0,0,94115
4221,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.3,19.3,0,50,0,16.36,5626,0,San Francisco,0,1,NA,37.744409999999995,-122.486764,0,19.3,0,0,Offer E,42959,0,0,0,0,1,2,0.0,16.36,0.0,19.3,0,0,94116
4222,1,0,0,0,45,1,0,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),112.2,5031.85,0,57,3,28.72,3091,0,San Francisco,1,1,DSL,37.770533,-122.445121,0,112.2,0,0,None,38756,1,0,0,1,45,0,151.0,1292.4,0.0,5031.85,0,0,94117
4223,1,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.3,220.4,0,35,27,9.74,4275,0,San Francisco,0,1,Cable,37.781304,-122.461522,0,70.3,0,0,None,38955,0,0,0,0,3,1,60.0,29.22,0.0,220.4,0,0,94118
4224,0,0,1,0,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.6,1416.5,0,46,0,37.83,4890,0,San Francisco,0,0,NA,37.776718,-122.49578100000001,1,19.6,0,2,None,42476,0,0,1,0,71,0,0.0,2685.93,0.0,1416.5,0,0,94121
4225,1,0,1,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,158.35,0,29,0,4.98,4964,0,San Francisco,0,1,NA,37.760412,-122.48496599999999,1,20.25,0,9,None,55504,0,0,1,0,8,2,0.0,39.84,0.0,158.35,1,0,94122
4226,0,0,1,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.85,256.6,1,61,32,44.34,4062,1,San Francisco,0,0,Cable,37.800253999999995,-122.436975,1,78.884,0,1,Offer E,22920,0,0,1,0,3,4,82.0,133.02,0.0,256.6,0,0,94123
4227,1,0,1,1,69,1,0,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),80.65,5542.55,0,48,53,40.36,4618,0,San Francisco,0,1,DSL,37.731505,-122.38453200000001,1,80.65,3,5,None,33177,1,0,1,1,69,1,2938.0,2784.84,0.0,5542.55,0,0,94124
4228,1,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,68.5,68.5,1,39,12,30.62,5753,1,San Francisco,0,1,DSL,37.736534999999996,-122.45732,1,71.24000000000002,0,1,Offer E,20643,0,0,1,0,1,0,0.0,30.62,0.0,68.5,0,0,94127
4229,0,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),115.75,8443.7,0,75,24,44.89,6205,0,San Francisco,1,0,DSL,37.797526,-122.46453100000001,1,115.75,0,2,Offer A,2240,1,0,1,0,72,0,2026.0,3232.08,0.0,8443.7,0,0,94129
4230,1,0,0,0,11,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,73.5,791.75,1,30,33,38.88,4509,1,San Francisco,0,1,DSL,37.820894,-122.369725,0,76.44,0,0,None,1458,0,0,0,0,11,5,261.0,427.68,0.0,791.75,0,0,94130
4231,1,0,0,0,71,1,1,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),80.6,5708.2,0,51,21,12.27,5447,0,San Francisco,1,1,Cable,37.746699,-122.44283300000001,0,80.6,0,0,None,27906,1,0,0,1,71,2,1199.0,871.17,0.0,5708.2,0,0,94131
4232,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.95,69.95,1,29,51,13.04,5341,1,San Francisco,0,0,Fiber Optic,37.722302,-122.491129,0,72.748,0,0,Offer E,26297,0,0,0,0,1,0,0.0,13.04,0.0,69.95,1,0,94132
4233,0,0,1,0,33,0,No phone service,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),59.55,2016.3,0,52,7,0.0,5980,0,San Francisco,1,0,Fiber Optic,37.802071000000005,-122.411004,1,59.55,0,7,Offer C,26831,1,0,1,1,33,0,141.0,0.0,0.0,2016.3,0,0,94133
4234,0,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.05,326.65,0,62,0,41.51,4336,0,San Francisco,0,0,NA,37.721052,-122.413573,0,19.05,0,0,Offer D,40137,0,0,0,0,16,1,0.0,664.16,0.0,326.65,0,0,94134
4235,0,1,1,0,56,1,1,Fiber optic,1,1,0,0,One year,0,Electronic check,95.65,5471.75,0,80,27,11.55,6335,0,Palo Alto,1,0,Fiber Optic,37.444314,-122.149996,1,95.65,0,10,Offer B,16198,1,0,1,0,56,2,1477.0,646.8000000000002,21.71,5471.75,0,0,94301
4236,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.95,19.95,0,58,0,38.84,2732,0,Palo Alto,0,0,NA,37.458090000000006,-122.115398,0,19.95,0,0,None,45499,0,0,0,0,1,2,0.0,38.84,0.0,19.95,0,0,94303
4237,1,0,0,0,5,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,70.05,346.4,1,52,29,14.26,4944,1,Palo Alto,1,1,DSL,37.386978000000006,-122.177746,0,72.852,0,0,None,1723,0,2,0,1,5,5,0.0,71.3,0.0,346.4,0,1,94304
4238,1,0,1,1,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.4,1061.6,0,45,0,41.56,4194,0,Stanford,0,1,NA,37.424341999999996,-122.165641,1,19.4,2,1,None,13386,0,0,1,0,57,0,0.0,2368.92,0.0,1061.6,0,0,94305
4239,1,0,1,1,56,0,No phone service,DSL,0,1,0,0,One year,1,Credit card (automatic),36.1,1971.5,0,61,28,0.0,5092,0,Palo Alto,1,1,Fiber Optic,37.416159,-122.13133700000002,1,36.1,1,1,None,24492,0,0,1,0,56,0,0.0,0.0,0.0,1971.5,0,1,94306
4240,1,0,0,0,8,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,94.0,773.65,1,59,15,23.89,2632,1,San Mateo,1,1,DSL,37.590421,-122.306467,0,97.76,0,0,None,32488,0,1,0,0,8,3,116.0,191.12,0.0,773.65,0,0,94401
4241,0,0,1,1,22,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,61.15,1422.05,1,21,33,42.98,4626,1,San Mateo,1,0,DSL,37.556634,-122.317723,1,63.596,3,1,Offer D,23393,0,0,1,0,22,0,0.0,945.56,0.0,1422.05,1,1,94402
4242,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.75,19.75,0,59,0,41.28,4099,0,San Mateo,0,0,NA,37.538309000000005,-122.305109,0,19.75,0,0,None,37926,0,1,0,0,1,1,0.0,41.28,0.0,19.75,0,0,94403
4243,0,0,0,1,40,1,0,DSL,1,0,1,0,Month-to-month,1,Credit card (automatic),64.1,2460.35,0,63,10,20.13,5056,0,San Mateo,0,0,Fiber Optic,37.556094,-122.27243700000001,0,64.1,1,0,None,31882,1,0,0,0,40,2,246.0,805.1999999999998,0.0,2460.35,0,0,94404
4244,1,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.75,856.5,0,62,0,7.67,2610,0,Alameda,0,1,NA,37.774633,-122.27443400000001,1,19.75,3,0,None,58555,0,0,0,0,46,1,0.0,352.82,0.0,856.5,0,0,94501
4245,1,0,1,1,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.7,1275.85,0,47,0,3.65,4235,0,Alameda,0,1,NA,37.724817,-122.22436299999998,1,19.7,1,0,None,13996,0,0,0,0,63,0,0.0,229.95,0.0,1275.85,0,0,94502
4246,1,0,1,1,68,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,110.2,7467.5,0,51,75,18.47,4108,0,Danville,1,1,Fiber Optic,37.791481,-121.903253,1,110.2,3,1,None,19777,0,0,1,1,68,0,5601.0,1255.96,0.0,7467.5,0,0,94506
4247,1,0,1,1,69,1,0,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),106.35,7261.75,0,38,24,42.9,6315,0,Alamo,0,1,Fiber Optic,37.855717,-121.994813,1,106.35,2,1,None,15187,1,0,1,1,69,0,1743.0,2960.1,0.0,7261.75,0,0,94507
4248,0,0,1,0,56,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,90.55,5116.6,0,63,20,2.8,6161,0,Angwin,1,0,Fiber Optic,38.542448,-122.419923,1,90.55,0,1,None,3641,1,0,1,0,56,0,0.0,156.79999999999995,0.0,5116.6,0,1,94508
4249,0,0,1,1,10,1,0,DSL,0,1,0,1,One year,1,Mailed check,65.9,660.05,0,32,14,42.0,5289,0,Antioch,1,0,DSL,37.980057,-121.801599,1,65.9,2,1,Offer D,90891,0,0,1,1,10,0,0.0,420.0,0.0,660.05,0,1,94509
4250,1,0,0,0,63,1,1,Fiber optic,1,1,1,0,One year,0,Credit card (automatic),104.5,6590.8,0,26,85,21.45,4908,0,Benicia,1,1,Cable,38.113533000000004,-122.11926000000001,0,104.5,0,0,None,25578,1,1,0,0,63,2,5602.0,1351.35,0.0,6590.8,1,0,94510
4251,0,0,1,1,24,0,No phone service,DSL,1,1,0,1,Two year,1,Mailed check,52.5,1208.15,0,34,75,0.0,3303,0,Bethel Island,1,0,Fiber Optic,38.050558,-121.646924,1,52.5,3,1,Offer C,2379,1,0,1,1,24,1,0.0,0.0,0.0,1208.15,0,1,94511
4252,0,0,0,0,19,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,56.1,1033.9,0,54,27,36.88,3367,0,Birds Landing,1,0,Cable,38.140719,-121.838298,0,56.1,0,0,Offer D,138,0,1,0,0,19,1,279.0,700.72,0.0,1033.9,0,0,94512
4253,1,0,1,1,22,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,88.75,1885.15,0,53,56,11.39,5585,0,Brentwood,1,1,Fiber Optic,37.908242,-121.682472,1,88.75,3,1,Offer D,26577,0,0,1,0,22,0,1056.0,250.58,0.0,1885.15,0,0,94513
4254,1,0,1,0,29,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,84.45,2467.1,1,37,13,28.37,2651,1,Byron,0,1,DSL,37.83323,-121.60146100000001,1,87.82799999999999,0,0,None,10153,0,0,0,0,29,2,0.0,822.73,0.0,2467.1,0,1,94514
4255,1,0,1,0,13,1,1,DSL,0,0,1,1,One year,1,Mailed check,75.3,989.45,1,20,90,41.22,4800,1,Calistoga,1,1,DSL,38.629618,-122.593216,1,78.312,0,1,Offer D,7384,0,3,1,1,13,4,891.0,535.86,0.0,989.45,1,0,94515
4256,0,0,1,0,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),26.0,2006.95,0,44,0,14.15,6170,0,Clayton,0,0,NA,37.881842,-121.84811100000002,1,26.0,0,1,None,14239,0,0,1,0,70,2,0.0,990.5,0.0,2006.95,0,0,94517
4257,0,0,1,0,49,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,99.4,5025,0,20,46,12.39,4725,0,Concord,1,0,Cable,37.950247999999995,-122.02245500000001,1,99.4,0,1,None,27394,0,0,1,1,49,1,0.0,607.11,0.0,5025.0,1,1,94518
4258,0,1,1,0,43,1,1,Fiber optic,1,0,1,1,One year,1,Mailed check,109.55,4830.25,1,74,14,8.75,5863,1,Concord,1,0,Cable,37.990118,-122.012188,1,113.932,0,7,Offer B,18650,1,0,1,0,43,3,67.62,376.25,0.0,4830.25,0,1,94519
4259,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.6,59.75,1,38,0,13.28,5000,1,Concord,0,0,NA,38.013825,-122.039144,0,19.6,0,0,Offer E,36186,0,1,0,0,3,3,0.0,39.84,0.0,59.75,0,0,94520
4260,1,0,1,1,42,1,0,DSL,0,0,1,1,One year,0,Electronic check,73.15,3088.25,0,54,23,14.8,2531,0,Concord,1,1,Fiber Optic,37.971421,-121.97150400000001,1,73.15,2,1,None,39888,1,0,1,1,42,2,710.0,621.6,0.0,3088.25,0,0,94521
4261,1,0,0,0,57,1,0,DSL,0,1,0,0,One year,1,Mailed check,54.65,3134.7,0,57,20,9.32,4223,0,Pleasant Hill,0,1,Fiber Optic,37.953379999999996,-122.07688600000002,0,54.65,0,0,None,32685,1,0,0,0,57,1,627.0,531.24,0.0,3134.7,0,0,94523
4262,1,1,0,0,2,1,0,DSL,1,0,1,0,Month-to-month,0,Bank transfer (automatic),66.4,94.55,1,73,26,5.57,4522,1,Crockett,1,1,Cable,38.049292,-122.22841499999998,0,69.05600000000001,0,0,None,3193,0,0,0,0,2,0,25.0,11.14,0.0,94.55,0,0,94525
4263,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),115.55,8312.4,0,23,59,1.67,5076,0,Danville,1,0,DSL,37.815459000000004,-121.977203,1,115.55,0,1,None,32873,1,0,1,1,72,0,490.43,120.24,0.0,8312.4,1,1,94526
4264,0,1,0,0,46,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.45,4863.85,0,65,30,41.17,4103,0,El Cerrito,1,0,DSL,37.924838,-122.28914499999999,0,104.45,0,0,Offer B,23141,0,0,0,1,46,1,0.0,1893.82,36.78,4863.85,0,1,94530
4265,1,1,1,0,66,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),100.05,6871.9,1,71,15,49.85,4512,1,Fairfield,0,1,Cable,38.287136,-122.02711000000001,1,104.052,0,6,None,77683,1,0,1,0,66,4,1031.0,3290.1,0.0,6871.9,0,0,94533
4266,1,0,0,0,62,1,1,Fiber optic,1,1,0,1,One year,0,Electronic check,102.0,6529.25,1,63,23,8.08,5090,1,Travis Afb,0,1,Cable,38.265899,-121.93946100000001,0,106.08,0,0,Offer B,9978,1,0,0,1,62,6,1502.0,500.96,0.0,6529.25,0,0,94535
4267,0,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),91.15,6637.9,0,53,26,2.95,4311,0,Fremont,1,0,DSL,37.572272999999996,-121.964583,1,91.15,0,4,None,66543,1,0,1,1,72,1,0.0,212.4,0.0,6637.9,0,1,94536
4268,1,0,1,1,35,1,0,Fiber optic,0,1,1,0,One year,1,Electronic check,89.7,3165.6,0,50,57,1.53,2775,0,Fremont,0,1,DSL,37.505767999999996,-121.96247199999999,1,89.7,3,5,Offer C,56126,1,0,1,0,35,0,0.0,53.55,0.0,3165.6,0,1,94538
4269,1,0,1,0,17,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Credit card (automatic),90.2,1454.15,1,62,10,12.06,2026,1,Fremont,1,1,DSL,37.516791,-121.89911699999999,1,93.80799999999999,0,1,Offer D,46917,0,2,1,0,17,1,145.0,205.02,0.0,1454.15,0,0,94539
4270,0,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Electronic check,92.4,6786.1,0,20,48,37.45,5527,0,Hayward,1,0,Fiber Optic,37.674002,-122.076796,1,92.4,0,8,None,60274,1,0,1,1,72,1,325.73,2696.4,0.0,6786.1,1,1,94541
4271,0,0,1,1,28,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.9,543,0,64,0,21.91,2987,0,Hayward,0,0,NA,37.656695,-122.04836100000001,1,19.9,1,9,Offer C,11147,0,0,1,0,28,0,0.0,613.48,0.0,543.0,0,0,94542
4272,1,0,1,0,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.15,1327.15,1,19,0,13.2,6484,1,Hayward,0,1,NA,37.639215,-122.037554,1,25.15,0,1,Offer B,72993,0,1,1,0,56,4,0.0,739.1999999999998,0.0,1327.15,1,0,94544
4273,0,0,0,0,31,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),79.85,2404.15,1,58,13,16.63,2554,1,Hayward,0,0,Cable,37.62984,-122.120843,0,83.044,0,0,None,27311,1,0,0,0,31,3,313.0,515.53,0.0,2404.15,0,0,94545
4274,1,0,0,0,45,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),18.85,867.3,0,47,0,40.59,2653,0,Castro Valley,0,1,NA,37.708327000000004,-122.083473,0,18.85,0,0,None,41698,0,0,0,0,45,2,0.0,1826.55,0.0,867.3,0,0,94546
4275,0,0,0,0,1,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,25.75,25.75,0,23,0,15.22,2569,0,Hercules,0,0,NA,37.991259,-122.214945,0,25.75,0,0,None,22479,0,0,0,0,1,0,0.0,15.22,0.0,25.75,1,0,94547
4276,0,0,0,0,2,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,49.6,114.7,1,26,29,21.28,3599,1,Lafayette,0,0,DSL,37.907777,-122.12716100000002,0,51.583999999999996,0,0,Offer E,23996,0,1,0,0,2,1,33.0,42.56,0.0,114.7,1,0,94549
4277,0,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.95,109.5,0,40,0,43.19,5554,0,Livermore,0,0,NA,37.571748,-121.65956200000001,0,20.95,0,0,None,75929,0,0,0,0,6,0,0.0,259.14,0.0,109.5,0,0,94550
4278,0,0,1,0,48,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,97.05,4692.95,0,29,59,47.64,5893,0,Castro Valley,1,0,Fiber Optic,37.722727,-122.02157,1,97.05,0,4,None,13212,0,0,1,1,48,1,0.0,2286.7200000000007,0.0,4692.95,1,1,94552
4279,1,0,1,1,25,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),25.4,546.85,0,61,0,19.56,5250,0,Martinez,0,1,NA,38.014457,-122.11543200000001,1,25.4,4,8,Offer C,46677,0,0,1,0,25,2,0.0,489.0,0.0,546.85,0,0,94553
4280,1,0,1,1,64,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.7,1274.05,0,28,0,14.93,5431,0,Fremont,0,1,NA,37.555473,-122.080312,1,19.7,1,3,Offer B,33883,0,0,1,0,64,0,0.0,955.52,0.0,1274.05,1,0,94555
4281,1,0,0,0,50,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Mailed check,35.0,1782.4,0,51,20,0.0,5629,0,Moraga,0,1,Fiber Optic,37.827946000000004,-122.10718500000002,0,35.0,0,0,Offer B,16510,0,0,0,0,50,0,0.0,0.0,0.0,1782.4,0,1,94556
4282,0,0,1,1,52,1,1,Fiber optic,0,0,1,1,One year,0,Bank transfer (automatic),101.25,5301.1,0,20,52,44.79,5954,0,Napa,1,0,Cable,38.489789,-122.27011,1,101.25,1,1,Offer B,63947,0,0,1,1,52,0,0.0,2329.08,0.0,5301.1,1,1,94558
4283,1,1,1,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.2,280.35,0,70,8,6.03,4444,0,Napa,0,1,Cable,38.232389000000005,-122.32494399999999,1,70.2,0,5,None,26894,0,0,1,0,4,1,0.0,24.12,30.75,280.35,0,1,94559
4284,0,1,0,0,32,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,90.95,2897.95,0,80,4,31.57,5936,0,Newark,0,0,Fiber Optic,37.504133,-122.032347,0,90.95,0,0,Offer C,42491,0,0,0,0,32,0,0.0,1010.24,25.55,2897.95,0,1,94560
4285,1,0,1,1,45,1,1,DSL,1,1,1,0,Two year,0,Credit card (automatic),73.85,3371,0,21,26,25.69,5264,0,Oakley,0,1,DSL,37.999406,-121.686241,1,73.85,1,9,Offer B,27607,1,1,1,0,45,1,0.0,1156.05,0.0,3371.0,1,1,94561
4286,1,0,1,0,9,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,88.05,801.3,0,49,21,22.41,2715,0,Orinda,0,1,DSL,37.873915999999994,-122.20522,1,88.05,0,3,None,17964,0,0,1,1,9,0,16.83,201.69,0.0,801.3,0,1,94563
4287,0,1,1,0,66,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),105.95,6975.25,1,68,12,27.75,6117,1,Pinole,1,0,Fiber Optic,37.996462,-122.29371599999999,1,110.18799999999999,0,1,None,16717,1,0,1,0,66,0,837.0,1831.5,0.0,6975.25,0,0,94564
4288,1,0,0,1,3,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,91.85,257.05,1,53,23,43.72,2704,1,Pittsburg,1,1,Cable,38.006046999999995,-121.91683400000001,0,95.524,0,0,None,78816,0,0,0,1,3,4,59.0,131.16,0.0,257.05,0,0,94565
4289,0,0,0,0,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.1,1079.45,0,45,0,26.25,5755,0,Pleasanton,0,0,NA,37.633361,-121.86239499999999,0,20.1,0,0,Offer B,36669,0,0,0,0,54,1,0.0,1417.5,0.0,1079.45,0,0,94566
4290,0,0,1,1,1,0,No phone service,DSL,0,0,1,0,Month-to-month,0,Electronic check,40.1,40.1,1,42,13,0.0,5434,1,Pope Valley,0,0,Fiber Optic,38.672708,-122.40321899999999,1,41.70399999999999,2,1,None,494,1,2,1,0,1,5,0.0,0.0,0.0,40.1,0,1,94567
4291,0,0,1,1,64,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),110.3,6997.3,0,49,23,21.16,5574,0,Dublin,0,0,Cable,37.713926,-121.928425,1,110.3,1,7,Offer B,29636,1,0,1,1,64,1,0.0,1354.24,0.0,6997.3,0,1,94568
4292,0,1,0,0,31,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.9,2217.15,1,70,2,15.43,2560,1,Port Costa,0,0,Cable,38.035707,-122.196821,0,76.85600000000002,0,0,None,173,0,0,0,0,31,4,44.0,478.33,0.0,2217.15,0,0,94569
4293,0,0,0,0,14,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,89.8,1129.1,1,57,32,10.3,4107,1,Rio Vista,0,0,Cable,38.148862,-121.737696,0,93.39200000000001,0,0,Offer D,5246,0,2,0,1,14,1,361.0,144.20000000000005,0.0,1129.1,0,0,94571
4294,0,0,0,0,12,1,0,Fiber optic,1,0,1,0,One year,1,Credit card (automatic),85.15,979.05,0,61,19,15.97,2452,0,Rodeo,0,0,DSL,38.027218,-122.23463000000001,0,85.15,0,0,Offer D,8506,0,2,0,0,12,1,0.0,191.64,0.0,979.05,0,1,94572
4295,1,1,1,0,67,1,0,DSL,1,1,0,0,One year,1,Bank transfer (automatic),60.95,4119.4,0,79,12,42.07,5792,0,Saint Helena,0,1,Fiber Optic,38.581354,-122.296283,1,60.95,0,7,Offer A,9423,1,0,1,0,67,2,0.0,2818.69,17.19,4119.4,0,1,94574
4296,0,0,1,1,35,1,1,DSL,1,0,1,0,Month-to-month,0,Electronic check,72.25,2568.55,1,28,90,25.27,5898,1,Deer Park,1,0,DSL,38.554383,-122.474773,1,75.14,2,1,None,223,1,0,1,0,35,3,2312.0,884.4499999999998,0.0,2568.55,1,0,94576
4297,0,0,0,0,45,1,1,DSL,1,0,0,1,Two year,0,Mailed check,73.55,3349.1,0,60,15,44.29,2280,0,San Leandro,0,0,Cable,37.717196,-122.15933799999999,0,73.55,0,0,Offer B,41871,1,0,0,1,45,0,0.0,1993.05,0.0,3349.1,0,1,94577
4298,1,0,0,0,10,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,46.0,492.1,0,45,14,13.51,3903,0,San Leandro,0,1,Cable,37.704384000000005,-122.126703,0,46.0,0,0,Offer D,36568,0,0,0,0,10,0,69.0,135.1,0.0,492.1,0,0,94578
4299,0,1,0,0,29,1,1,DSL,1,1,0,0,Month-to-month,1,Bank transfer (automatic),58.55,1718.95,0,68,22,8.88,2044,0,San Leandro,0,0,Fiber Optic,37.687264,-122.15728,0,58.55,0,0,Offer C,19815,0,0,0,0,29,1,0.0,257.52000000000004,33.1,1718.95,0,1,94579
4300,0,0,0,0,24,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),24.6,605.25,0,58,0,42.66,4147,0,San Lorenzo,0,0,NA,37.676249,-122.132415,0,24.6,0,0,Offer C,26240,0,0,0,0,24,0,0.0,1023.84,0.0,605.25,0,0,94580
4301,1,0,1,1,66,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.75,1344.5,0,62,0,31.53,4485,0,San Ramon,0,1,NA,37.766556,-121.97678400000001,1,19.75,2,7,None,44078,0,0,1,0,66,0,0.0,2080.98,0.0,1344.5,0,0,94583
4302,1,0,0,0,51,1,0,Fiber optic,1,0,1,0,One year,0,Mailed check,86.35,4267.15,0,51,13,27.3,5311,0,Suisun City,0,1,DSL,38.197907,-122.01725800000001,0,86.35,0,0,Offer B,39279,0,0,0,0,51,3,555.0,1392.3,0.0,4267.15,0,0,94585
4303,0,0,1,0,45,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.5,1121.05,0,35,0,42.32,3146,0,Sunol,0,0,NA,37.587494,-121.86285600000001,1,25.5,0,6,Offer B,790,0,0,1,0,45,1,0.0,1904.4,0.0,1121.05,0,0,94586
4304,0,0,1,0,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.0,918.7,0,54,0,13.13,4066,0,Union City,0,0,NA,37.59485,-122.051521,1,19.0,0,3,Offer B,66472,0,0,1,0,49,2,0.0,643.37,0.0,918.7,0,0,94587
4305,0,0,1,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.55,521.8,0,44,0,49.96,5758,0,Pleasanton,0,0,NA,37.685052,-121.91206100000001,1,19.55,0,6,Offer C,28568,0,0,1,0,29,1,0.0,1448.84,0.0,521.8,0,0,94588
4306,1,0,1,1,40,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),110.1,4469.1,0,59,22,11.5,2283,0,Vallejo,0,1,Fiber Optic,38.161321,-122.271588,1,110.1,3,6,Offer B,42209,1,0,1,1,40,3,0.0,460.0,0.0,4469.1,0,1,94589
4307,0,1,0,0,37,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.55,3580.3,1,66,2,3.3,4448,1,Vallejo,0,0,Cable,38.104704999999996,-122.24738700000002,0,100.412,0,0,None,37218,0,1,0,0,37,5,0.0,122.1,0.0,3580.3,0,1,94590
4308,1,0,0,0,25,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.75,1729.35,0,42,18,40.11,3080,0,Vallejo,0,1,Cable,38.105733,-122.18633799999999,0,69.75,0,0,Offer C,51665,0,0,0,0,25,0,31.13,1002.75,0.0,1729.35,0,1,94591
4309,0,0,0,0,22,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,50.6,1073.3,0,34,8,0.0,2854,0,Vallejo,1,0,DSL,38.093701,-122.27658899999999,0,50.6,0,0,None,159,0,0,0,1,22,1,0.0,0.0,0.0,1073.3,0,1,94592
4310,1,0,0,0,72,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),65.6,4566.5,0,36,9,0.0,4369,0,Walnut Creek,1,1,Fiber Optic,37.862128000000006,-122.075197,0,65.6,0,0,None,18024,1,0,0,1,72,4,411.0,0.0,0.0,4566.5,0,0,94595
4311,0,0,0,0,7,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Credit card (automatic),40.1,293.3,1,36,21,0.0,4414,1,Walnut Creek,0,0,Cable,37.900662,-122.05278200000001,0,41.70399999999999,0,0,None,40917,0,0,0,1,7,0,6.16,0.0,0.0,293.3,0,1,94596
4312,1,0,1,1,33,1,0,DSL,0,1,1,1,Two year,0,Credit card (automatic),82.1,2603.1,0,44,30,1.62,2281,0,Walnut Creek,1,1,Fiber Optic,37.916647999999995,-122.00848300000001,1,82.1,1,1,Offer C,26022,1,0,1,1,33,0,781.0,53.46,0.0,2603.1,0,0,94598
4313,0,0,0,0,23,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,79.1,1783.75,0,22,46,15.18,3619,0,Yountville,0,0,Fiber Optic,38.421458,-122.365048,0,79.1,0,0,None,2873,1,0,0,0,23,0,0.0,349.14,0.0,1783.75,1,1,94599
4314,1,1,0,0,24,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.25,2440.15,1,65,33,28.98,4287,1,Oakland,0,1,Cable,37.776523,-122.219268,0,105.3,0,0,None,54876,0,1,0,1,24,2,805.0,695.52,0.0,2440.15,0,0,94601
4315,0,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,79.55,79.55,1,58,16,32.13,5082,1,Oakland,0,0,Fiber Optic,37.803883,-122.208417,0,82.73200000000001,0,0,None,28900,0,0,0,0,1,1,0.0,32.13,0.0,79.55,0,0,94602
4316,1,0,0,0,69,1,1,DSL,1,1,1,1,Two year,0,Mailed check,90.65,6322.1,0,42,22,47.43,6487,0,Oakland,1,1,DSL,37.739113,-122.175602,0,90.65,0,0,None,31392,1,0,0,1,69,3,1391.0,3272.67,0.0,6322.1,0,0,94603
4317,0,0,0,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.55,57.4,0,37,0,11.27,2774,0,Oakland,0,0,NA,37.758019,-122.138678,0,20.55,2,0,None,42854,0,0,0,0,3,2,0.0,33.81,0.0,57.4,0,0,94605
4318,1,0,0,0,56,1,0,DSL,0,1,1,1,One year,1,Bank transfer (automatic),75.75,4284.65,0,61,13,18.42,6487,0,Oakland,0,1,Fiber Optic,37.792489,-122.24431399999999,0,75.75,0,0,Offer B,41876,1,0,0,1,56,2,0.0,1031.52,0.0,4284.65,0,1,94606
4319,1,0,0,0,65,1,1,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),110.0,7138.65,0,61,10,33.11,6351,0,Oakland,1,1,Fiber Optic,37.80707,-122.29740100000001,0,110.0,0,0,None,21054,1,0,0,1,65,0,714.0,2152.15,0.0,7138.65,0,0,94607
4320,1,0,1,0,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,20.85,1539.75,0,55,0,44.82,4837,0,Emeryville,0,1,NA,37.83726,-122.287648,1,20.85,0,5,None,24589,0,0,1,0,71,4,0.0,3182.22,0.0,1539.75,0,0,94608
4321,0,1,0,0,14,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),80.35,1058.1,0,73,3,7.34,3276,0,Oakland,1,0,DSL,37.834340999999995,-122.26437,0,80.35,0,0,None,21097,0,0,0,0,14,2,32.0,102.76,32.71,1058.1,0,0,94609
4322,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.15,123.8,0,57,10,33.75,4840,0,Oakland,0,0,Fiber Optic,37.808731,-122.238708,0,70.15,0,0,None,29964,0,1,0,0,2,1,12.0,67.5,0.0,123.8,0,0,94610
4323,0,0,0,0,32,1,1,Fiber optic,0,0,1,0,One year,0,Electronic check,84.05,2781.85,1,44,15,40.26,3553,1,Oakland,0,0,DSL,37.828416,-122.21600500000001,0,87.412,0,0,None,36517,0,2,0,0,32,2,0.0,1288.32,0.0,2781.85,0,1,94611
4324,1,0,0,0,40,1,0,DSL,1,0,0,1,Month-to-month,0,Electronic check,67.45,2731,0,28,58,39.05,4714,0,Oakland,1,1,DSL,37.809014000000005,-122.26973899999999,0,67.45,0,0,None,11702,0,0,0,1,40,1,158.4,1562.0,0.0,2731.0,1,1,94612
4325,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.75,20.75,0,49,0,36.28,2791,0,Oakland,0,1,NA,37.84551,-122.23518100000001,0,20.75,0,0,None,15438,0,0,0,0,1,2,0.0,36.28,0.0,20.75,0,0,94618
4326,1,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.1,89.1,1,44,3,16.06,2905,1,Oakland,0,1,DSL,37.787186,-122.14633,0,92.664,0,0,None,24518,0,0,0,1,1,6,0.0,16.06,0.0,89.1,0,0,94619
4327,0,0,0,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.9,497.3,0,25,42,30.99,4562,0,Oakland,0,0,Fiber Optic,37.750553000000004,-122.197175,0,69.9,0,0,None,30751,0,0,0,0,7,4,0.0,216.93,0.0,497.3,1,1,94621
4328,0,0,1,0,15,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,51.1,711.15,0,60,5,31.13,4858,0,Berkeley,0,0,DSL,37.866009000000005,-122.28622800000001,1,51.1,0,1,None,15638,0,2,1,0,15,1,0.0,466.95,0.0,711.15,0,1,94702
4329,0,0,1,1,17,1,1,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,94.4,1607.2,1,57,13,25.79,4103,1,Berkeley,1,0,Cable,37.863843,-122.27568400000001,1,98.17600000000002,0,1,Offer D,19763,0,1,1,0,17,1,209.0,438.43,0.0,1607.2,0,0,94703
4330,1,0,0,0,19,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,78.25,1490.95,1,59,28,20.26,3666,1,Berkeley,1,1,Fiber Optic,37.871415999999996,-122.246597,0,81.38000000000002,0,0,Offer D,21205,0,2,0,0,19,3,0.0,384.94000000000005,0.0,1490.95,0,1,94704
4331,1,0,0,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.55,1898.1,0,43,0,39.08,6305,0,Berkeley,0,1,NA,37.858897999999996,-122.24051200000001,0,25.55,0,0,None,12448,0,0,0,0,71,2,0.0,2774.68,0.0,1898.1,0,0,94705
4332,0,0,1,1,54,1,1,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),60.0,3273.95,0,22,73,8.53,4798,0,Albany,0,0,DSL,37.890274,-122.29519199999999,1,60.0,3,6,None,15882,1,0,1,0,54,2,2390.0,460.62,0.0,3273.95,1,0,94706
4333,1,0,1,0,31,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),90.55,2929.75,0,47,21,22.42,5722,0,Berkeley,0,1,Cable,37.897753,-122.27939099999999,1,90.55,0,4,Offer C,11889,1,0,1,0,31,1,615.0,695.0200000000002,0.0,2929.75,0,0,94707
4334,0,0,0,0,11,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,76.4,838.7,0,46,20,36.52,4033,0,Berkeley,0,0,Cable,37.897743,-122.263124,0,76.4,0,0,None,10737,0,0,0,0,11,2,168.0,401.72,0.0,838.7,0,0,94708
4335,0,1,0,0,18,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.95,1443.65,0,70,23,25.7,3878,0,Berkeley,1,0,Cable,37.878554,-122.26608999999999,0,84.95,0,0,None,10147,0,0,0,0,18,0,332.0,462.6,4.76,1443.65,0,0,94709
4336,0,1,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),110.1,7746.7,0,77,23,14.12,5232,0,Berkeley,0,0,DSL,37.872902,-122.30370800000001,0,110.1,0,0,Offer A,8157,1,0,0,0,72,0,0.0,1016.64,44.81,7746.7,0,1,94710
4337,0,1,0,0,71,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),99.65,6951.15,0,73,13,34.36,4241,0,Richmond,0,0,Cable,37.945288,-122.383941,0,99.65,0,0,Offer A,28450,0,0,0,0,71,1,904.0,2439.56,3.33,6951.15,0,0,94801
4338,1,1,0,0,5,0,No phone service,DSL,0,0,1,0,Month-to-month,0,Credit card (automatic),45.4,214.75,0,74,4,0.0,2599,0,El Sobrante,1,1,Fiber Optic,37.963995000000004,-122.288296,0,45.4,0,0,None,25399,1,0,0,0,5,0,0.0,0.0,0.0,214.75,0,1,94803
4339,1,0,1,0,38,1,1,DSL,0,0,0,1,One year,0,Credit card (automatic),69.0,2669.45,0,34,16,32.11,4487,0,Richmond,1,1,Fiber Optic,37.921034000000006,-122.341798,1,69.0,0,2,Offer C,39089,1,0,1,1,38,1,427.0,1220.18,0.0,2669.45,0,0,94804
4340,1,0,0,1,5,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),48.65,235.2,0,57,21,13.54,3307,0,Richmond,0,1,DSL,37.941456,-122.320968,0,48.65,2,0,None,13984,1,2,0,0,5,1,0.0,67.69999999999999,0.0,235.2,0,1,94805
4341,1,1,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.15,92.65,1,78,28,43.66,5655,1,San Pablo,0,1,Fiber Optic,37.980269,-122.34263500000002,0,45.916000000000004,0,0,None,55720,0,1,0,0,2,5,26.0,87.32,0.0,92.65,0,0,94806
4342,0,1,0,0,52,1,1,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),59.85,3103.25,0,78,3,34.0,5085,0,San Rafael,1,0,Fiber Optic,37.972662,-122.491452,0,59.85,0,0,Offer B,40239,0,0,0,0,52,1,0.0,1768.0,19.16,3103.25,0,1,94901
4343,0,1,0,0,8,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.75,606.25,1,74,7,13.8,4174,1,San Rafael,0,0,DSL,38.018065,-122.546024,0,78.78,0,0,None,28403,0,1,0,0,8,3,42.0,110.4,0.0,606.25,0,0,94903
4344,0,0,0,0,68,1,1,DSL,0,1,1,1,Two year,1,Electronic check,80.65,5330.2,0,52,13,20.3,5914,0,Greenbrae,1,0,Cable,37.946616999999996,-122.563571,0,80.65,0,0,None,12010,0,0,0,1,68,1,0.0,1380.4,0.0,5330.2,0,1,94904
4345,1,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.55,1403.1,0,23,0,26.44,5366,0,Belvedere Tiburon,0,1,NA,37.885628999999994,-122.46858,1,20.55,2,8,Offer A,13065,0,0,1,0,69,2,0.0,1824.36,0.0,1403.1,1,0,94920
4346,0,0,1,0,42,1,1,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),66.4,2727.8,0,56,30,36.35,3773,0,Bodega,0,0,Cable,38.343282,-122.9755,1,66.4,0,4,None,584,1,0,1,0,42,0,0.0,1526.7,0.0,2727.8,0,1,94922
4347,0,0,0,0,50,1,0,Fiber optic,0,1,1,1,Two year,1,Mailed check,100.2,5038.45,0,36,9,15.1,5419,0,Bodega Bay,0,0,Fiber Optic,38.377165000000005,-123.037957,0,100.2,0,0,None,1785,1,0,0,1,50,0,0.0,755.0,0.0,5038.45,0,1,94923
4348,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.1,19.1,1,35,0,34.79,5890,1,Bolinas,0,0,NA,37.943087,-122.72379,0,19.1,0,0,None,1573,0,0,0,0,1,4,0.0,34.79,0.0,19.1,0,0,94924
4349,1,1,1,0,1,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,80.3,80.3,1,78,23,17.51,4138,1,Corte Madera,0,1,Cable,37.924014,-122.51169399999999,1,83.512,0,1,None,9038,0,2,1,0,1,2,0.0,17.51,0.0,80.3,0,0,94925
4350,1,0,1,0,33,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),44.55,1462.6,0,23,51,48.49,2422,0,Rohnert Park,0,1,Fiber Optic,38.347190000000005,-122.697822,1,44.55,0,6,Offer C,42544,0,0,1,0,33,1,746.0,1600.17,0.0,1462.6,1,0,94928
4351,0,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,150.6,0,43,0,41.57,3098,0,Dillon Beach,0,0,NA,38.24458,-122.956268,0,20.35,0,0,Offer E,330,0,0,0,0,7,1,0.0,290.99,0.0,150.6,0,0,94929
4352,1,0,1,1,64,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,91.8,5960.5,0,21,27,34.58,5371,0,Fairfax,1,1,Cable,37.971751,-122.611873,1,91.8,1,0,None,8486,0,0,0,0,64,1,1609.0,2213.12,0.0,5960.5,1,0,94930
4353,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.9,74.9,1,26,33,35.25,5919,1,Cotati,1,0,Fiber Optic,38.326215000000005,-122.71874199999999,0,77.89600000000002,0,0,None,7936,0,2,0,0,1,1,0.0,35.25,0.0,74.9,1,0,94931
4354,1,0,0,0,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.2,1192.3,0,47,0,47.17,5216,0,Forest Knolls,0,1,NA,38.010092,-122.68944199999999,0,20.2,0,0,None,1025,0,0,0,0,59,0,0.0,2783.03,0.0,1192.3,0,0,94933
4355,0,0,1,0,6,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,50.35,314.55,0,30,85,42.66,3442,0,Inverness,0,0,Fiber Optic,38.099323,-122.945723,1,50.35,0,10,Offer E,1004,0,0,1,0,6,0,267.0,255.96,0.0,314.55,0,0,94937
4356,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,18.8,56,0,44,0,6.61,3010,0,Lagunitas,0,0,NA,38.021772,-122.691744,0,18.8,0,0,Offer E,821,0,0,0,0,3,0,0.0,19.83,0.0,56.0,0,0,94938
4357,0,0,1,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.45,330.8,0,21,0,12.41,5184,0,Larkspur,0,0,NA,37.937082000000004,-122.53236899999999,1,20.45,0,3,None,6773,0,0,1,0,15,0,0.0,186.15,0.0,330.8,1,0,94939
4358,1,0,1,1,13,1,0,DSL,0,0,1,1,One year,1,Electronic check,64.75,877.35,0,59,21,13.32,4741,0,Marshall,0,1,Fiber Optic,38.129308,-122.83481499999999,1,64.75,1,1,None,406,0,0,1,1,13,0,184.0,173.16,0.0,877.35,0,0,94940
4359,0,0,0,0,23,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),98.7,2249.1,0,40,19,14.45,5781,0,Mill Valley,0,0,Fiber Optic,37.901371000000005,-122.572024,0,98.7,0,0,None,28727,0,0,0,1,23,2,0.0,332.35,0.0,2249.1,0,1,94941
4360,1,1,1,0,31,1,1,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,89.45,2807.65,0,76,18,46.06,5597,0,Novato,0,1,DSL,38.135897,-122.56368300000001,1,89.45,0,5,Offer C,16429,0,0,1,0,31,2,50.54,1427.86,31.58,2807.65,0,1,94945
4361,1,0,0,0,29,1,0,DSL,1,1,0,0,One year,1,Electronic check,58.75,1696.2,0,35,9,8.0,5198,0,Nicasio,0,1,Fiber Optic,38.065359,-122.665566,0,58.75,0,0,Offer C,607,1,0,0,0,29,1,153.0,232.0,0.0,1696.2,0,0,94946
4362,0,0,1,0,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.7,1032.05,0,62,0,29.18,4074,0,Novato,0,0,NA,38.112165999999995,-122.63438400000001,1,20.7,0,0,None,24741,0,0,0,0,49,2,0.0,1429.82,0.0,1032.05,0,0,94947
4363,0,0,1,0,56,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),85.6,4902.8,0,25,51,42.81,6483,0,Novato,0,0,DSL,38.067204,-122.524004,1,85.6,0,9,None,13361,0,0,1,0,56,0,250.04,2397.36,0.0,4902.8,1,1,94949
4364,0,0,0,0,63,1,1,DSL,1,1,0,1,Two year,1,Credit card (automatic),80.3,4995.35,0,50,26,31.34,5554,0,Olema,1,0,DSL,38.052209000000005,-122.775567,0,80.3,0,0,None,248,1,0,0,1,63,0,129.88,1974.42,0.0,4995.35,0,1,94950
4365,1,0,1,0,63,1,1,DSL,0,0,1,1,Two year,0,Credit card (automatic),79.8,5034.05,0,51,20,10.07,4073,0,Penngrove,1,1,DSL,38.325599,-122.642352,1,79.8,0,5,None,3777,1,0,1,1,63,2,0.0,634.41,0.0,5034.05,0,1,94951
4366,1,1,1,1,24,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,79.85,1857.75,0,66,28,4.06,3412,0,Petaluma,0,1,Fiber Optic,38.237018,-122.77871999999999,1,79.85,2,6,Offer C,31930,0,0,1,0,24,0,520.0,97.44,0.0,1857.75,0,0,94952
4367,1,1,1,0,36,1,0,DSL,0,0,0,0,One year,0,Credit card (automatic),54.1,1992.85,0,65,28,47.16,4017,0,Petaluma,1,1,Fiber Optic,38.235021,-122.557332,1,54.1,0,9,Offer C,35419,1,0,1,0,36,0,0.0,1697.7599999999998,1.09,1992.85,0,1,94954
4368,0,1,0,0,9,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.85,751.65,1,79,2,43.34,5242,1,Point Reyes Station,0,0,Fiber Optic,38.060264000000004,-122.830646,0,84.084,0,0,None,1885,0,0,0,0,9,7,15.0,390.06000000000006,0.0,751.65,0,0,94956
4369,1,0,0,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,24.75,66.95,1,36,20,0.0,3503,1,San Anselmo,0,1,DSL,37.99272,-122.575026,0,25.74,0,0,None,16849,0,0,0,0,3,4,13.0,0.0,0.0,66.95,0,0,94960
4370,0,0,1,0,21,1,0,DSL,1,0,1,1,One year,0,Mailed check,80.9,1714.95,0,55,19,11.27,5733,0,San Geronimo,1,0,Fiber Optic,38.004740000000005,-122.66371699999999,1,80.9,0,7,None,548,1,0,1,1,21,0,326.0,236.67,0.0,1714.95,0,0,94963
4371,1,0,1,1,13,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),24.5,343.6,0,31,0,48.7,5077,0,San Quentin,0,1,NA,37.942551,-122.491642,1,24.5,2,8,None,6448,0,0,1,0,13,0,0.0,633.1,0.0,343.6,0,0,94964
4372,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.15,20.15,0,25,0,18.63,3960,0,Sausalito,0,1,NA,37.848641,-122.51569199999999,1,20.15,2,7,Offer E,11213,0,0,1,0,1,0,0.0,18.63,0.0,20.15,1,0,94965
4373,0,0,1,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.05,520.1,0,52,0,13.06,2010,0,Stinson Beach,0,0,NA,37.921137,-122.65756200000001,1,20.05,2,7,Offer C,781,0,0,1,0,25,0,0.0,326.5,0.0,520.1,0,0,94970
4374,1,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.6,1387.45,0,64,0,16.13,6444,0,Tomales,0,1,NA,38.240769,-122.90104099999999,1,19.6,3,6,Offer A,384,0,0,1,0,71,1,0.0,1145.23,0.0,1387.45,0,0,94971
4375,1,0,0,0,66,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),114.3,7383.7,0,27,73,4.32,5303,0,Valley Ford,1,1,Fiber Optic,38.339996,-122.935056,0,114.3,0,0,Offer A,66,1,0,0,1,66,0,0.0,285.12,0.0,7383.7,1,1,94972
4376,0,0,0,0,45,1,0,Fiber optic,1,1,1,1,One year,1,Electronic check,100.3,4483.95,0,27,47,1.03,4868,0,Woodacre,0,0,Fiber Optic,38.005839,-122.638155,0,100.3,0,0,None,1449,0,0,0,1,45,0,210.75,46.35,0.0,4483.95,1,1,94973
4377,0,0,1,0,22,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),80.0,1706.45,0,20,41,45.1,2640,0,Alviso,0,0,DSL,37.449537,-121.994813,1,80.0,0,1,None,2147,0,0,1,0,22,1,0.0,992.2,0.0,1706.45,1,1,95002
4378,0,0,1,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),20.85,1327.4,0,57,0,7.91,5972,0,Aptos,0,0,NA,37.013471,-121.877877,1,20.85,0,5,Offer A,24227,0,0,1,0,67,0,0.0,529.97,0.0,1327.4,0,0,95003
4379,0,0,1,0,68,1,1,Fiber optic,0,0,1,0,Two year,1,Bank transfer (automatic),89.95,5974.3,0,30,82,28.36,5672,0,Aromas,1,0,DSL,36.878364000000005,-121.62978100000001,1,89.95,0,5,Offer A,3373,0,0,1,0,68,0,0.0,1928.48,0.0,5974.3,0,1,95004
4380,0,0,1,1,0,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.0, ,0,23,0,20.05,3763,0,Ben Lomond,0,0,NA,37.078873,-122.09038600000001,1,20.0,3,4,Offer E,6407,0,0,1,0,10,1,0.0,200.5,0.0,200.0,1,0,95005
4381,0,1,0,0,49,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),90.85,4515.85,1,76,16,44.88,5651,1,Boulder Creek,1,0,Cable,37.171727000000004,-122.14296100000001,0,94.484,0,0,Offer B,10520,0,0,0,0,49,5,723.0,2199.120000000001,0.0,4515.85,0,0,95006
4382,0,1,0,0,4,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,48.75,179.85,0,65,15,31.13,3048,0,Brookdale,0,0,DSL,37.106902000000005,-122.10000600000001,0,48.75,0,0,None,1007,0,0,0,0,4,1,0.0,124.52,0.0,179.85,0,1,95007
4383,1,0,1,0,63,1,1,DSL,1,1,0,1,One year,0,Credit card (automatic),80.0,5040.2,0,34,18,34.02,5540,0,Campbell,1,1,Cable,37.279689000000005,-121.954567,1,80.0,0,9,None,44976,1,0,1,1,63,1,907.0,2143.26,0.0,5040.2,0,0,95008
4384,0,0,1,0,2,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),79.7,165,1,25,29,28.86,3039,1,Capitola,1,0,DSL,36.977025,-121.95286399999999,1,82.88799999999999,0,1,None,9673,0,3,1,0,2,2,48.0,57.72,0.0,165.0,1,0,95010
4385,1,0,0,0,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.35,422.7,0,31,0,22.53,3721,0,Castroville,0,1,NA,36.784481,-121.759054,0,20.35,0,0,None,8582,0,0,0,0,21,1,0.0,473.13,0.0,422.7,0,0,95012
4386,1,0,1,1,55,1,0,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),57.55,3046.4,1,28,53,8.8,5463,1,Cupertino,0,1,Fiber Optic,37.306612,-122.080621,1,59.852,0,1,Offer B,54431,1,0,1,0,55,0,1615.0,484.00000000000006,0.0,3046.4,1,0,95014
4387,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.25,20.25,0,21,0,47.25,2448,0,Davenport,0,1,NA,37.114335,-122.23716200000001,0,20.25,2,0,Offer E,857,0,0,0,0,1,1,0.0,47.25,0.0,20.25,1,0,95017
4388,0,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.4,358.05,0,58,0,30.07,3561,0,Felton,0,0,NA,37.089110999999995,-122.06221299999999,0,19.4,0,0,Offer D,8728,0,0,0,0,17,0,0.0,511.19,0.0,358.05,0,0,95018
4389,1,0,0,0,30,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),100.4,2936.25,0,45,19,17.26,3778,0,Freedom,0,1,DSL,36.936228,-121.785559,0,100.4,0,0,Offer C,4753,0,0,0,1,30,1,0.0,517.8000000000002,0.0,2936.25,0,1,95019
4390,1,0,1,1,22,1,0,DSL,1,1,0,0,Month-to-month,1,Mailed check,57.95,1271.8,0,21,82,42.58,5036,0,Gilroy,0,1,Cable,37.03889,-121.52895500000001,1,57.95,3,9,Offer D,49968,1,0,1,1,22,1,1043.0,936.76,0.0,1271.8,1,0,95020
4391,0,0,0,0,9,1,0,DSL,0,0,1,0,Month-to-month,1,Bank transfer (automatic),59.5,530.05,0,33,20,39.19,4011,0,Escondido,0,0,DSL,33.141265000000004,-116.967221,0,59.5,0,0,Offer E,48690,1,0,0,0,9,0,0.0,352.71,0.0,530.05,0,1,92027
4392,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.2,19.2,0,57,0,32.78,3007,0,Los Gatos,0,1,NA,37.222842,-121.988727,1,19.2,3,10,None,13290,0,0,1,0,1,0,0.0,32.78,0.0,19.2,0,0,95030
4393,0,0,1,0,21,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.5,1808.7,1,50,32,42.22,2036,1,Los Gatos,0,0,Fiber Optic,37.233034,-121.947427,1,89.96000000000002,0,3,Offer D,24443,0,0,1,1,21,4,579.0,886.62,0.0,1808.7,0,0,95032
4394,1,0,0,0,19,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,59.55,1144.6,0,40,18,11.85,3949,0,Los Gatos,1,1,DSL,37.160194,-121.94561100000001,0,59.55,0,0,Offer D,10172,1,0,0,0,19,0,0.0,225.15,0.0,1144.6,0,1,95033
4395,0,0,1,1,69,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,103.95,7446.9,1,42,30,37.2,4283,1,Milpitas,1,0,Cable,37.441931,-121.878502,1,108.10799999999999,0,1,None,62848,0,0,1,1,69,4,2234.0,2566.8,0.0,7446.9,0,0,95035
4396,1,1,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,25.1,25.1,1,67,10,0.0,5437,1,Morgan Hill,0,1,Cable,37.161544,-121.649371,0,26.104000000000006,0,0,None,41707,0,0,0,0,1,0,0.0,0.0,0.0,25.1,0,1,95037
4397,0,0,1,0,72,1,1,Fiber optic,1,1,1,0,Two year,1,Bank transfer (automatic),103.95,7556.9,0,33,8,44.27,5096,0,Moss Landing,1,0,Fiber Optic,36.863303,-121.781632,1,103.95,0,10,Offer A,899,1,0,1,0,72,0,0.0,3187.44,0.0,7556.9,0,1,95039
4398,1,0,1,1,70,1,1,DSL,1,0,1,0,Two year,0,Credit card (automatic),68.95,4858.7,0,49,29,22.67,4858,0,Mount Hermon,1,1,DSL,37.051165999999995,-122.05619399999999,1,68.95,1,9,Offer A,77,0,2,1,0,70,2,1409.0,1586.9,0.0,4858.7,0,0,95041
4399,0,0,0,0,66,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Bank transfer (automatic),103.1,6595,0,33,20,43.14,6183,0,Paicines,1,0,DSL,36.525703,-120.952122,0,103.1,0,0,Offer A,813,1,0,0,1,66,2,131.9,2847.24,0.0,6595.0,0,1,95043
4400,0,0,1,1,7,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.7,149.05,0,20,76,0.0,3872,0,San Juan Bautista,0,0,Cable,36.810567999999996,-121.503022,1,24.7,2,3,None,3402,0,0,1,1,7,3,0.0,0.0,0.0,149.05,1,1,95045
4401,0,1,1,1,46,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,110.2,4972.1,0,76,16,20.42,4162,0,San Martin,0,0,Cable,37.084697,-121.606417,1,110.2,1,7,Offer B,5671,1,0,1,0,46,0,0.0,939.32,0.0,4972.1,0,1,95046
4402,1,0,0,0,39,0,No phone service,DSL,1,1,1,0,Month-to-month,1,Credit card (automatic),48.95,1880.85,1,27,53,0.0,3080,1,Santa Clara,0,1,Cable,37.351214,-121.952417,0,50.908,0,0,None,36349,1,0,0,0,39,3,0.0,0.0,0.0,1880.85,1,1,95050
4403,0,0,1,1,32,1,1,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),62.45,2045.55,0,29,51,33.28,5442,0,Santa Clara,1,0,DSL,37.348129,-121.98468999999999,1,62.45,1,9,Offer C,52986,0,0,1,1,32,0,0.0,1064.96,0.0,2045.55,1,1,95051
4404,1,0,0,0,24,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.55,2187.15,0,21,59,27.91,2007,0,Santa Clara,1,1,Fiber Optic,37.393553999999995,-121.96511399999999,0,89.55,0,0,None,13031,0,0,0,1,24,1,129.04,669.84,0.0,2187.15,1,1,95054
4405,1,0,1,1,6,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),83.55,477.55,1,47,7,26.91,4242,1,Santa Cruz,0,1,DSL,36.993451,-122.098858,1,86.89200000000001,0,1,None,43192,0,2,1,1,6,3,33.0,161.46,0.0,477.55,0,0,95060
4406,0,0,0,0,37,1,1,DSL,1,1,1,0,Month-to-month,1,Credit card (automatic),78.9,2976.95,0,43,4,42.41,3801,0,Santa Cruz,1,0,Fiber Optic,36.974575,-121.991149,0,78.9,0,0,None,36631,1,0,0,0,37,0,0.0,1569.1699999999996,0.0,2976.95,0,1,95062
4407,1,0,0,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,178.7,0,61,0,14.37,4577,0,Santa Cruz,0,1,NA,37.007882,-122.065975,0,20.35,1,0,None,4563,0,0,0,0,8,0,0.0,114.96,0.0,178.7,0,0,95064
4408,0,0,1,1,72,1,1,DSL,1,0,1,0,Two year,1,Bank transfer (automatic),71.45,5025.85,0,26,73,38.99,5656,0,Santa Cruz,1,0,DSL,37.031403999999995,-121.98186499999998,1,71.45,1,8,Offer A,8365,0,0,1,1,72,0,3669.0,2807.28,0.0,5025.85,1,0,95065
4409,1,1,1,0,71,0,No phone service,DSL,1,1,0,0,Two year,0,Credit card (automatic),46.35,3353.4,0,74,19,0.0,5421,0,Scotts Valley,1,1,Fiber Optic,37.070177,-122.010077,1,46.35,0,9,Offer A,14574,1,0,1,0,71,0,0.0,0.0,18.64,3353.4,0,1,95066
4410,0,0,1,0,16,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),94.65,1461.15,0,56,2,10.5,3050,0,Saratoga,0,0,Fiber Optic,37.257771999999996,-122.051824,1,94.65,0,3,Offer D,30589,0,0,1,1,16,0,0.0,168.0,0.0,1461.15,0,1,95070
4411,0,0,1,0,57,0,No phone service,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),49.9,2782.4,0,44,14,0.0,5866,0,Soquel,1,0,Cable,37.023669,-121.94646100000001,1,49.9,0,2,None,9823,1,2,1,1,57,1,0.0,0.0,0.0,2782.4,0,1,95073
4412,1,0,0,0,66,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),25.45,1699.15,0,40,0,32.22,4163,0,Watsonville,0,1,NA,36.931653999999995,-121.75238300000001,0,25.45,0,0,Offer A,81141,0,0,0,0,66,0,0.0,2126.52,0.0,1699.15,0,0,95076
4413,0,1,0,0,17,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.15,1496.9,1,80,31,30.37,5082,1,San Jose,1,0,DSL,37.34667,-121.91001899999999,0,92.716,0,0,Offer D,18197,0,1,0,0,17,6,464.0,516.29,0.0,1496.9,0,0,95110
4414,0,0,0,1,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.75,452.2,0,38,0,8.68,2143,0,San Jose,0,0,NA,37.284265000000005,-121.827673,0,20.75,2,0,Offer D,57748,0,0,0,0,21,0,0.0,182.28,0.0,452.2,0,0,95111
4415,1,0,1,0,66,1,1,DSL,1,1,0,0,Two year,1,Credit card (automatic),66.1,4428.45,0,43,15,37.71,5933,0,San Jose,1,1,Cable,37.343827000000005,-121.883119,1,66.1,0,9,Offer A,52334,0,1,1,0,66,3,66.43,2488.86,0.0,4428.45,0,1,95112
4416,0,0,1,0,17,1,1,DSL,0,1,1,1,Month-to-month,1,Bank transfer (automatic),75.4,1322.55,0,29,52,7.6,4852,0,San Jose,0,0,Cable,37.333851,-121.891147,1,75.4,0,5,Offer D,561,0,0,1,1,17,0,688.0,129.2,0.0,1322.55,1,0,95113
4417,1,0,0,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.45,70.45,1,42,9,42.87,3525,1,San Jose,0,1,Cable,37.350284,-121.852855,0,73.268,0,0,None,51706,0,4,0,0,1,3,0.0,42.87,0.0,70.45,0,0,95116
4418,1,0,1,0,58,1,0,DSL,1,1,0,0,One year,0,Credit card (automatic),60.3,3563.8,1,31,23,17.22,4026,1,San Jose,1,1,Cable,37.311088,-121.961786,1,62.712,0,1,Offer B,29914,0,0,1,0,58,0,820.0,998.76,0.0,3563.8,0,0,95117
4419,0,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),21.05,139.75,0,54,0,43.05,2158,0,San Jose,0,0,NA,37.255479,-121.88983799999998,1,21.05,3,5,None,31926,0,0,1,0,8,2,0.0,344.4,0.0,139.75,0,0,95118
4420,1,0,0,0,27,1,0,DSL,1,0,1,0,One year,0,Credit card (automatic),69.35,1927.3,0,19,26,36.39,2450,0,San Jose,1,1,Cable,37.233226,-121.78809,0,69.35,0,0,None,10155,1,0,0,1,27,1,501.0,982.53,0.0,1927.3,1,0,95119
4421,1,0,1,0,34,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Mailed check,88.85,3000.25,0,28,48,13.97,4014,0,San Jose,0,1,Cable,37.186141,-121.843554,1,88.85,0,10,None,37090,0,0,1,1,34,0,0.0,474.98,0.0,3000.25,1,1,95120
4422,1,0,0,0,30,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),97.0,3021.3,0,44,16,12.17,4126,0,San Jose,0,1,Fiber Optic,37.304681,-121.809955,0,97.0,0,0,None,37127,0,0,0,1,30,1,483.0,365.1,0.0,3021.3,0,0,95121
4423,1,0,0,0,33,1,0,DSL,0,1,1,0,Month-to-month,1,Credit card (automatic),66.4,2245.4,0,19,51,45.72,3843,0,San Jose,1,1,Fiber Optic,37.32886,-121.83456699999999,0,66.4,0,0,None,59841,0,0,0,1,33,0,0.0,1508.76,0.0,2245.4,1,1,95122
4424,1,0,0,1,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,24.75,24.75,1,56,63,0.0,3001,1,San Jose,0,1,Fiber Optic,37.238758000000004,-121.828375,0,25.74,3,0,None,59632,0,3,0,0,1,4,0.0,0.0,0.0,24.75,0,0,95123
4425,1,0,1,1,14,1,1,DSL,1,1,0,1,Month-to-month,0,Mailed check,69.2,944.65,0,52,76,2.96,2871,0,San Jose,0,1,DSL,37.257063,-121.92303700000001,1,69.2,3,8,Offer D,45257,0,0,1,1,14,4,0.0,41.44,0.0,944.65,0,1,95124
4426,0,0,0,1,16,1,1,Fiber optic,0,0,0,0,One year,1,Credit card (automatic),79.5,1264.2,0,30,69,27.23,5040,0,San Jose,0,0,Cable,37.294926000000004,-121.89476299999998,0,79.5,3,0,Offer D,46185,1,1,0,0,16,2,87.23,435.68,0.0,1264.2,0,1,95125
4427,0,0,0,0,49,1,0,Fiber optic,0,0,1,1,Two year,0,Credit card (automatic),100.65,4917.75,0,49,27,11.11,5499,0,San Jose,1,0,Fiber Optic,37.327069,-121.91681899999999,0,100.65,0,0,None,27023,1,0,0,1,49,0,1328.0,544.39,0.0,4917.75,0,0,95126
4428,1,0,1,1,19,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,103.3,2012.7,1,34,24,28.04,2349,1,San Jose,1,1,Fiber Optic,37.375156,-121.79586699999999,1,107.432,0,1,Offer D,60620,1,2,1,1,19,2,483.0,532.76,0.0,2012.7,0,0,95127
4429,0,0,1,1,70,1,1,DSL,1,1,1,0,Two year,0,Bank transfer (automatic),79.7,5743.3,0,44,19,8.36,4848,0,San Jose,1,0,Fiber Optic,37.316146,-121.93628500000001,1,79.7,1,3,Offer A,32804,1,1,1,0,70,2,1091.0,585.1999999999998,0.0,5743.3,0,0,95128
4430,0,0,1,1,32,1,0,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),61.4,1864.65,0,49,17,46.66,2649,0,San Jose,0,0,DSL,37.305622,-122.000887,1,61.4,1,3,None,37570,1,0,1,0,32,1,31.7,1493.12,0.0,1864.65,0,1,95129
4431,0,0,0,0,18,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.8,1221.65,0,35,20,34.12,2421,0,San Jose,0,0,Cable,37.277592,-121.98647700000001,0,69.8,0,0,Offer D,13481,0,0,0,0,18,0,244.0,614.16,0.0,1221.65,0,0,95130
4432,1,0,0,0,37,0,No phone service,DSL,1,1,0,0,Two year,1,Mailed check,40.55,1390.85,0,26,69,0.0,4050,0,San Jose,0,1,Fiber Optic,37.387027,-121.897775,0,40.55,0,0,None,26389,1,0,0,1,37,0,0.0,0.0,0.0,1390.85,1,1,95131
4433,0,0,0,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.65,302.35,0,36,22,23.5,5396,0,San Jose,0,0,DSL,37.424655,-121.74841,0,75.65,0,0,None,40568,0,0,0,0,4,0,0.0,94.0,0.0,302.35,0,1,95132
4434,0,0,1,0,16,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Electronic check,90.7,1374.9,0,19,52,27.83,4839,0,San Jose,1,0,DSL,37.371862,-121.860349,1,90.7,0,2,Offer D,26032,0,1,1,1,16,1,715.0,445.28,0.0,1374.9,1,0,95133
4435,1,0,1,0,17,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.5,1336.9,0,31,8,46.71,3591,0,San Jose,0,1,Fiber Optic,37.42765,-121.945416,1,80.5,0,7,Offer D,9657,0,0,1,0,17,1,0.0,794.07,0.0,1336.9,0,1,95134
4436,0,0,0,1,19,1,0,DSL,1,1,0,0,Month-to-month,1,Electronic check,60.6,1297.8,0,52,20,36.48,2463,0,San Jose,1,0,Cable,37.28682,-121.723877,0,60.6,3,0,Offer D,15798,0,0,0,0,19,1,0.0,693.1199999999999,0.0,1297.8,0,1,95135
4437,1,0,1,0,60,1,1,Fiber optic,0,0,1,1,Two year,0,Credit card (automatic),101.15,6067.4,0,27,48,10.05,5301,0,San Jose,1,1,Fiber Optic,37.270938,-121.851046,1,101.15,0,0,None,36944,0,0,0,1,60,0,2912.0,603.0,0.0,6067.4,1,0,95136
4438,1,0,1,1,51,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.95,1222.25,0,46,0,16.85,5461,0,San Jose,0,1,NA,37.246064000000004,-121.749494,1,24.95,2,7,None,14792,0,1,1,0,51,1,0.0,859.35,0.0,1222.25,0,0,95138
4439,1,0,1,1,28,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.3,487.95,0,30,0,19.18,2948,0,San Jose,0,1,NA,37.218705,-121.762429,1,20.3,2,8,None,7023,0,0,1,0,28,0,0.0,537.04,0.0,487.95,0,0,95139
4440,1,0,0,0,43,1,0,DSL,0,1,0,1,Two year,1,Electronic check,60.0,2548.55,0,64,13,21.64,4614,0,Mount Hamilton,0,1,Fiber Optic,37.382909000000005,-121.634151,0,60.0,0,0,None,38,0,0,0,1,43,0,331.0,930.52,0.0,2548.55,0,0,95140
4441,1,0,1,0,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,20.25,835.5,0,49,0,45.75,5940,0,San Jose,0,1,NA,37.339533,-121.777179,1,20.25,0,10,None,44103,0,0,1,0,42,2,0.0,1921.5,0.0,835.5,0,0,95148
4442,1,0,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,78.5,242.05,1,39,8,31.88,3567,1,Stockton,0,1,Cable,37.959706,-121.287669,0,81.64,0,0,None,7071,0,1,0,0,3,1,0.0,95.64,0.0,242.05,0,1,95202
4443,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.75,44.75,0,35,21,40.87,4118,0,Stockton,0,0,Fiber Optic,37.954089,-121.329761,0,44.75,0,0,None,16357,0,0,0,0,1,2,0.0,40.87,0.0,44.75,0,1,95203
4444,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,63.75,1,24,0,25.75,3398,1,Stockton,0,0,NA,37.974498,-121.31956799999999,0,19.85,0,0,Offer E,30476,0,0,0,0,3,6,0.0,77.25,0.0,63.75,1,0,95204
4445,0,0,0,0,63,1,1,Fiber optic,1,1,1,0,Two year,0,Credit card (automatic),98.0,6218.45,0,49,21,23.62,5989,0,Stockton,1,0,DSL,37.965695000000004,-121.260051,0,98.0,0,0,None,34138,0,0,0,0,63,1,1306.0,1488.0600000000004,0.0,6218.45,0,0,95205
4446,1,1,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.9,260.9,1,77,3,2.98,4367,1,Stockton,0,1,Fiber Optic,37.902421999999994,-121.44002900000001,0,83.096,0,0,None,49657,0,0,0,0,3,1,8.0,8.94,0.0,260.9,0,0,95206
4447,1,0,1,0,68,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,107.7,7320.9,0,25,48,24.01,5015,0,Stockton,0,1,Fiber Optic,38.002125,-121.324979,1,107.7,0,2,Offer A,49965,1,1,1,1,68,1,0.0,1632.68,0.0,7320.9,1,1,95207
4448,0,1,0,0,30,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.7,2967.35,1,73,9,43.61,3548,1,Stockton,0,0,DSL,38.044523,-121.34804799999999,0,103.68799999999999,0,0,None,30814,0,2,0,0,30,2,267.0,1308.3,0.0,2967.35,0,0,95209
4449,0,0,0,0,60,1,1,Fiber optic,0,1,1,1,Two year,0,Electronic check,104.7,6333.8,0,23,51,35.47,6186,0,Stockton,1,0,Cable,38.033219,-121.29743300000001,0,104.7,0,0,None,40611,0,0,0,1,60,1,323.02,2128.2,0.0,6333.8,1,1,95210
4450,1,0,0,0,15,1,1,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),58.6,939.7,1,29,65,14.79,2003,1,Stockton,0,1,Cable,38.049457000000004,-121.21653,0,60.943999999999996,0,0,Offer D,6951,1,1,0,0,15,3,611.0,221.85,0.0,939.7,1,0,95212
4451,1,1,0,0,45,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),93.9,4200.25,0,76,18,15.65,3960,0,Stockton,0,1,Fiber Optic,37.946282000000004,-121.139499,0,93.9,0,0,Offer B,23789,0,0,0,0,45,0,756.0,704.25,0.0,4200.25,0,0,95215
4452,0,0,1,0,70,1,0,DSL,1,1,1,1,Two year,0,Credit card (automatic),86.45,5950.2,0,31,5,31.15,5950,0,Stockton,1,0,Fiber Optic,38.029728999999996,-121.387999,1,86.45,0,0,Offer A,19109,1,0,0,1,70,0,298.0,2180.5,0.0,5950.2,0,0,95219
4453,1,0,1,0,10,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.5,1037.75,1,35,20,1.09,4501,1,Acampo,1,1,Fiber Optic,38.200231,-121.23503400000001,1,102.44,0,1,Offer D,6317,0,0,1,1,10,4,208.0,10.9,0.0,1037.75,0,0,95220
4454,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.4,93.4,0,26,0,22.54,4402,0,Angels Camp,0,1,NA,38.071327000000004,-120.632221,0,19.4,0,0,None,4264,0,0,0,0,4,0,0.0,90.16,0.0,93.4,1,0,95222
4455,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.45,50.45,1,39,19,23.7,2806,1,Arnold,1,0,Fiber Optic,38.321529999999996,-120.23635800000001,0,52.468,0,0,Offer E,5159,0,3,0,0,1,4,0.0,23.7,0.0,50.45,0,0,95223
4456,0,0,1,0,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.95,1614.9,0,38,0,26.64,6146,0,Avery,0,0,NA,38.208335999999996,-120.33993799999999,1,24.95,0,2,Offer A,115,0,0,1,0,68,0,0.0,1811.52,0.0,1614.9,0,0,95224
4457,1,0,1,1,22,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Bank transfer (automatic),75.0,1573.95,0,50,19,38.82,4040,0,Burson,0,1,DSL,38.183918,-120.898817,1,75.0,2,1,Offer D,27,0,0,1,0,22,4,0.0,854.04,0.0,1573.95,0,1,95225
4458,1,0,1,1,38,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,94.65,3624.3,1,25,33,49.7,3498,1,Campo Seco,1,1,Cable,38.233878999999995,-120.86166599999999,1,98.436,0,1,None,75,0,1,1,0,38,4,1196.0,1888.6,0.0,3624.3,1,0,95226
4459,0,0,0,0,1,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),100.25,100.25,1,45,19,20.23,5797,1,Clements,0,0,Fiber Optic,38.227284999999995,-121.02788999999999,0,104.26,0,0,Offer E,722,0,0,0,1,1,3,0.0,20.23,0.0,100.25,0,0,95227
4460,1,0,1,0,18,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,78.2,1468.75,0,55,19,31.79,2831,0,Copperopolis,1,1,DSL,37.943954,-120.67108,1,78.2,0,6,Offer D,2633,1,2,1,0,18,1,0.0,572.22,0.0,1468.75,0,1,95228
4461,1,0,0,0,29,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.2,2607.6,0,50,17,2.05,4561,0,Farmington,0,1,Fiber Optic,37.956963,-120.863055,0,94.2,0,0,None,596,1,0,0,1,29,1,443.0,59.45,0.0,2607.6,0,0,95230
4462,0,0,0,0,16,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,88.45,1422.1,1,44,6,17.8,5186,1,French Camp,1,0,Fiber Optic,37.873283,-121.29203400000002,0,91.988,0,0,Offer D,5094,0,1,0,1,16,1,85.0,284.8,0.0,1422.1,0,0,95231
4463,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.85,69.85,1,51,21,12.13,4548,1,Glencoe,0,1,Cable,38.358464,-120.57930400000001,0,72.64399999999998,0,0,Offer E,21,0,1,0,0,1,4,0.0,12.13,0.0,69.85,0,0,95232
4464,1,0,0,0,12,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Bank transfer (automatic),81.7,858.6,1,44,3,18.38,2850,1,Hathaway Pines,1,1,Cable,38.184914,-120.364085,0,84.96799999999999,0,0,Offer D,335,0,2,0,0,12,4,0.0,220.56,0.0,858.6,0,1,95233
4465,1,0,0,0,31,0,No phone service,DSL,0,0,1,1,One year,1,Electronic check,50.05,1523.4,0,35,5,0.0,4529,0,Linden,1,1,Fiber Optic,38.047746000000004,-121.030499,0,50.05,0,0,None,3148,0,0,0,1,31,1,0.0,0.0,0.0,1523.4,0,1,95236
4466,1,0,0,0,4,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.9,324.3,1,27,51,43.06,4669,1,Lockeford,0,1,DSL,38.166790999999996,-121.14206999999999,0,83.096,0,0,Offer E,3205,0,2,0,1,4,3,0.0,172.24,0.0,324.3,1,1,95237
4467,0,0,1,0,48,1,1,DSL,0,0,0,1,One year,1,Mailed check,69.55,3435.6,0,45,15,17.03,2478,0,Lodi,1,0,Fiber Optic,38.123544,-121.15907800000001,1,69.55,0,3,None,45755,1,0,1,1,48,0,515.0,817.44,0.0,3435.6,0,0,95240
4468,0,0,0,0,15,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),25.4,399.6,1,22,0,45.84,2853,1,Lodi,0,0,NA,38.128087,-121.4078,0,25.4,0,0,Offer D,22073,0,0,0,0,15,4,0.0,687.6,0.0,399.6,1,0,95242
4469,1,0,0,0,50,1,0,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),90.1,4549.45,0,34,22,15.37,6435,0,Mokelumne Hill,1,1,DSL,38.304194,-120.592431,0,90.1,0,0,None,2718,1,0,0,0,50,0,1001.0,768.5,0.0,4549.45,0,0,95245
4470,1,0,0,0,7,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),44.65,322.5,0,22,46,26.76,4300,0,Mountain Ranch,0,1,Fiber Optic,38.264262,-120.515133,0,44.65,0,0,None,1692,0,0,0,0,7,0,148.0,187.32,0.0,322.5,1,0,95246
4471,1,1,1,0,41,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),83.75,3273.55,1,74,20,45.84,4995,1,Murphys,1,1,Cable,38.147852,-120.440124,1,87.10000000000002,0,1,Offer B,4353,0,0,1,0,41,2,655.0,1879.44,0.0,3273.55,0,0,95247
4472,1,0,1,1,68,1,0,Fiber optic,1,0,0,0,Two year,0,Credit card (automatic),80.35,5375.15,0,25,41,24.08,5954,0,San Andreas,1,1,Cable,38.196496999999994,-120.61688999999998,1,80.35,3,8,Offer A,3930,0,0,1,0,68,0,2204.0,1637.4399999999996,0.0,5375.15,1,0,95249
4473,0,1,1,0,26,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),98.1,2510.7,0,79,11,18.66,3114,0,Sheep Ranch,1,0,Cable,38.244806,-120.417301,1,98.1,0,8,Offer C,88,0,1,1,0,26,1,276.0,485.16,44.17,2510.7,0,0,95250
4474,1,0,0,0,57,0,No phone service,DSL,0,0,1,1,Two year,0,Credit card (automatic),53.35,3090.05,0,33,28,0.0,5461,0,Vallecito,1,1,Fiber Optic,38.055562,-120.456298,0,53.35,0,0,None,460,1,0,0,1,57,0,865.0,0.0,0.0,3090.05,0,0,95251
4475,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.55,61.05,0,60,0,40.98,3889,0,Valley Springs,0,0,NA,38.156971,-120.849231,0,19.55,0,0,None,11266,0,0,0,0,3,2,0.0,122.94,0.0,61.05,0,0,95252
4476,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.9,20.9,1,21,0,15.73,5421,1,Wallace,0,0,NA,38.192608,-120.957842,0,20.9,0,0,Offer E,304,0,0,0,0,1,1,0.0,15.73,0.0,20.9,1,0,95254
4477,1,0,1,1,19,1,0,DSL,1,0,0,0,One year,1,Bank transfer (automatic),48.95,955.6,0,59,21,11.75,2394,0,West Point,0,1,Cable,38.41935,-120.469545,1,48.95,1,1,Offer D,2198,0,0,1,0,19,0,0.0,223.25,0.0,955.6,0,1,95255
4478,0,0,0,0,3,1,0,DSL,0,0,1,0,Month-to-month,1,Electronic check,54.2,140.4,0,50,5,41.38,3167,0,Wilseyville,0,0,Cable,38.392686,-120.415951,0,54.2,0,0,None,435,0,0,0,0,3,0,7.0,124.14,0.0,140.4,0,0,95257
4479,0,0,0,0,59,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,24.45,1493.1,0,64,0,41.23,6196,0,Woodbridge,0,0,NA,38.169605,-121.31096399999998,0,24.45,0,0,Offer B,4176,0,0,0,0,59,0,0.0,2432.57,0.0,1493.1,0,0,95258
4480,0,0,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.4,69.4,1,47,13,33.46,2404,1,Atwater,0,0,Fiber Optic,37.321233,-120.65635400000001,1,72.176,0,1,Offer E,27808,0,1,1,0,1,2,0.0,33.46,0.0,69.4,0,0,95301
4481,1,0,1,0,42,0,No phone service,DSL,1,0,1,0,Month-to-month,1,Bank transfer (automatic),40.15,1626.05,0,37,7,0.0,4348,0,Ballico,0,1,Fiber Optic,37.4695,-120.672724,1,40.15,0,1,Offer B,809,0,0,1,0,42,2,0.0,0.0,0.0,1626.05,0,1,95303
4482,0,0,0,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.9,541.15,1,62,28,46.79,5159,1,Big Oak Flat,0,0,DSL,37.818589,-120.25699499999999,0,77.89600000000002,0,0,Offer E,167,0,4,0,0,7,3,152.0,327.53,0.0,541.15,0,0,95305
4483,1,0,1,0,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.6,1784.9,0,58,0,11.74,4879,0,Catheys Valley,0,1,NA,37.394411,-120.12726200000002,1,25.6,0,1,Offer A,986,0,0,1,0,67,0,0.0,786.58,0.0,1784.9,0,0,95306
4484,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.35,70.35,0,63,27,14.42,2722,0,Ceres,0,1,Cable,37.553469,-120.952825,0,70.35,0,0,None,32881,0,0,0,0,1,0,0.0,14.42,0.0,70.35,0,0,95307
4485,1,0,1,0,66,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),91.7,6075.9,0,19,58,23.27,5453,0,Columbia,1,1,Cable,38.085839,-120.37855,1,91.7,0,1,Offer A,2144,1,0,1,1,66,0,0.0,1535.82,0.0,6075.9,1,1,95310
4486,0,0,0,0,61,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Mailed check,89.2,5500.6,0,60,27,14.52,5536,0,Coulterville,1,0,DSL,37.722127,-120.110174,0,89.2,0,0,Offer B,2271,0,0,0,1,61,0,0.0,885.72,0.0,5500.6,0,1,95311
4487,1,0,1,1,4,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),24.1,73.1,0,55,0,16.68,4463,0,Cressey,0,1,NA,37.420273,-120.66526999999999,1,24.1,2,1,Offer E,55,0,0,1,0,4,0,0.0,66.72,0.0,73.1,0,0,95312
4488,0,1,1,0,42,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),74.15,3229.4,1,76,23,2.9,2322,1,Crows Landing,0,0,Fiber Optic,37.435664,-121.04905600000001,1,77.11600000000001,0,1,Offer B,1508,0,0,1,0,42,5,0.0,121.8,0.0,3229.4,0,1,95313
4489,0,0,1,1,64,1,1,DSL,0,1,0,0,One year,1,Bank transfer (automatic),53.85,3399.85,0,53,25,17.07,4954,0,Delhi,0,0,DSL,37.422961,-120.76549299999999,1,53.85,2,10,Offer B,10159,0,0,1,0,64,0,0.0,1092.48,0.0,3399.85,0,1,95315
4490,0,1,1,0,54,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),115.6,6431.05,0,79,12,43.71,4337,0,Denair,1,0,Fiber Optic,37.524721,-120.757977,1,115.6,0,2,Offer B,5513,1,0,1,0,54,1,772.0,2360.34,0.0,6431.05,0,0,95316
4491,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.75,19.75,0,58,0,1.61,5809,0,El Nido,0,1,NA,37.127386,-120.506422,0,19.75,0,0,Offer E,808,0,1,0,0,1,1,0.0,1.61,0.0,19.75,0,0,95317
4492,1,0,1,1,54,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.05,1230.9,0,19,0,41.58,4039,0,El Portal,0,1,NA,37.654551,-119.822984,1,24.05,2,7,Offer B,579,0,0,1,0,54,2,0.0,2245.32,0.0,1230.9,1,0,95318
4493,0,0,0,1,18,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.3,454.65,0,45,0,30.22,3416,0,Escalon,0,0,NA,37.818543,-121.00690700000001,0,25.3,2,0,Offer D,11474,0,0,0,0,18,1,0.0,543.96,0.0,454.65,0,0,95320
4494,1,0,0,0,3,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,84.3,235.05,0,46,26,13.72,5828,0,Groveland,0,1,Fiber Optic,37.902968,-119.66754399999999,0,84.3,0,0,Offer E,3680,0,0,0,1,3,1,61.0,41.16,0.0,235.05,0,0,95321
4495,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.1,70.1,1,58,33,46.17,2007,1,Gustine,0,0,DSL,37.147197999999996,-121.12016100000001,0,72.904,0,0,Offer E,7872,0,0,0,0,1,1,0.0,46.17,0.0,70.1,0,1,95322
4496,0,0,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.75,6595.9,0,41,20,15.58,5096,0,Hickman,1,0,Fiber Optic,37.605926000000004,-120.69955,1,89.75,1,1,Offer A,1055,1,0,1,1,72,1,1319.0,1121.76,0.0,6595.9,0,0,95323
4497,1,1,1,0,60,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,97.95,5867,0,76,21,17.05,6150,0,Hilmar,1,1,Fiber Optic,37.394535999999995,-120.89074699999999,1,97.95,0,10,Offer B,7177,0,0,1,0,60,0,0.0,1023.0,0.0,5867.0,0,1,95324
4498,0,0,1,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.0,196.35,0,37,0,49.19,5837,0,Hornitos,0,0,NA,37.479926,-120.230424,1,20.0,1,8,Offer D,128,0,0,1,0,11,3,0.0,541.0899999999998,0.0,196.35,0,0,95325
4499,0,0,0,1,12,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,78.3,909.25,1,34,28,35.8,3545,1,Hughson,0,0,DSL,37.5923,-120.85328799999999,0,81.432,0,0,Offer D,6822,0,0,0,0,12,3,255.0,429.6,0.0,909.25,0,0,95326
4500,1,0,1,1,61,1,0,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),103.9,6449.15,0,37,19,43.08,4079,0,Jamestown,1,1,Cable,37.84771,-120.486589,1,103.9,1,3,Offer B,9559,1,0,1,1,61,0,0.0,2627.88,0.0,6449.15,0,1,95327
4501,0,0,0,0,39,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.7,762.45,0,23,0,29.79,3733,0,Keyes,0,0,NA,37.555631,-120.911653,0,20.7,0,0,None,2130,0,0,0,0,39,3,0.0,1161.81,0.0,762.45,1,0,95328
4502,1,0,0,0,55,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.8,5283.95,1,40,32,47.38,4089,1,La Grange,0,1,Cable,37.666587,-120.41151699999999,0,100.67200000000001,0,0,Offer B,1749,0,0,0,1,55,5,1691.0,2605.9,0.0,5283.95,0,0,95329
4503,0,0,0,0,17,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,94.4,1617.5,1,57,25,21.82,2825,1,Lathrop,0,0,Fiber Optic,37.808209999999995,-121.308401,0,98.17600000000002,0,0,Offer D,10834,0,0,0,0,17,5,404.0,370.94,0.0,1617.5,0,0,95330
4504,1,0,0,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.15,785.75,0,36,0,34.37,4422,0,Le Grand,0,1,NA,37.249377,-120.249581,0,20.15,0,0,None,3256,0,1,0,0,37,2,0.0,1271.6899999999996,0.0,785.75,0,0,95333
4505,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,26.0,1776,0,60,0,26.98,5374,0,Livingston,0,0,NA,37.361987,-120.74839399999999,1,26.0,0,8,Offer A,12672,0,0,1,0,72,0,0.0,1942.56,0.0,1776.0,0,0,95334
4506,1,1,1,0,72,1,1,DSL,0,1,1,0,Two year,0,Credit card (automatic),77.35,5396.25,0,73,10,33.68,6202,0,Long Barn,1,1,Fiber Optic,38.109125,-120.078597,1,77.35,0,4,Offer A,683,1,0,1,0,72,0,540.0,2424.96,0.0,5396.25,0,0,95335
4507,0,0,0,0,8,1,0,DSL,1,0,0,1,Month-to-month,0,Bank transfer (automatic),66.05,574.5,0,34,14,33.54,4157,0,Manteca,0,0,Fiber Optic,37.830267,-121.20101799999999,0,66.05,0,0,Offer E,36738,1,0,0,1,8,0,0.0,268.32,0.0,574.5,0,1,95336
4508,0,0,1,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,400.3,0,27,0,49.51,5657,0,Manteca,0,0,NA,37.750822,-121.238423,1,19.9,2,2,Offer D,19867,0,0,1,0,22,2,0.0,1089.22,0.0,400.3,1,0,95337
4509,0,0,0,0,1,1,0,Fiber optic,0,1,1,0,Month-to-month,0,Electronic check,84.3,84.3,1,27,65,1.63,2172,1,Mariposa,0,0,Fiber Optic,37.526790999999996,-119.99436999999999,0,87.67200000000001,0,0,None,10226,0,0,0,0,1,2,0.0,1.63,0.0,84.3,1,0,95338
4510,0,0,0,0,38,1,1,DSL,0,1,0,1,Month-to-month,0,Credit card (automatic),68.15,2656.3,0,61,24,21.19,3371,0,Merced,0,0,DSL,37.255637,-120.49353700000002,0,68.15,0,0,None,59289,1,0,0,1,38,1,63.75,805.22,0.0,2656.3,0,1,95340
4511,1,0,0,1,17,1,0,DSL,0,1,1,1,One year,0,Electronic check,80.85,1445.95,0,25,73,45.92,3913,0,Midpines,1,1,DSL,37.581496,-119.97276200000002,0,80.85,1,0,None,433,1,0,0,1,17,0,1056.0,780.64,0.0,1445.95,1,0,95345
4512,0,1,0,0,70,1,1,DSL,0,1,1,0,Two year,1,Bank transfer (automatic),75.5,5212.65,0,79,3,47.27,6024,0,Mi Wuk Village,1,0,Cable,38.121601,-120.13391499999999,0,75.5,0,0,Offer A,1278,1,0,0,0,70,0,15.64,3308.9,0.0,5212.65,0,1,95346
4513,0,1,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),92.45,6440.25,1,78,7,25.77,5697,1,Merced,1,0,DSL,37.40122,-120.514191,1,96.148,0,0,None,23100,1,0,0,0,72,1,0.0,1855.44,0.0,6440.25,0,1,95348
4514,0,0,0,0,28,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.6,2244.95,0,62,5,33.84,2951,0,Modesto,0,0,DSL,37.671806,-121.007575,0,80.6,0,0,None,52872,0,0,0,1,28,0,112.0,947.52,0.0,2244.95,0,0,95350
4515,0,0,0,0,15,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),83.2,1130,0,60,29,10.43,4096,0,Modesto,0,0,Fiber Optic,37.621458000000004,-121.012295,0,83.2,0,0,None,47536,0,0,0,0,15,1,328.0,156.45,0.0,1130.0,0,0,95351
4516,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),87.55,6463.15,0,59,53,44.61,5341,0,Modesto,1,1,Fiber Optic,37.639029,-120.964772,1,87.55,3,1,None,27135,1,0,1,1,72,1,0.0,3211.92,0.0,6463.15,0,1,95354
4517,0,1,1,0,11,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.55,1131.2,1,78,15,1.28,3172,1,Modesto,1,0,Cable,37.672906,-120.94659399999999,1,103.53200000000001,0,1,Offer D,47613,0,0,1,0,11,2,170.0,14.08,0.0,1131.2,0,0,95355
4518,1,1,0,0,8,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,81.25,585.95,1,66,29,5.02,3812,1,Modesto,1,1,Cable,37.716186,-121.02583600000001,0,84.5,0,0,None,26055,0,1,0,0,8,4,170.0,40.16,0.0,585.95,0,0,95356
4519,0,0,1,0,57,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),109.4,6252.7,0,20,73,8.01,6026,0,Modesto,1,0,Fiber Optic,37.670526,-120.877572,1,109.4,0,10,Offer B,13343,1,1,1,1,57,1,0.0,456.57,0.0,6252.7,1,1,95357
4520,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.95,19.95,1,52,0,8.03,4860,1,Modesto,0,1,NA,37.612612,-121.10856799999999,1,19.95,3,1,None,30668,0,0,1,0,1,1,0.0,8.03,0.0,19.95,0,0,95358
4521,0,0,1,0,46,0,No phone service,DSL,1,1,1,0,Month-to-month,0,Electronic check,45.55,2062.15,0,50,30,0.0,5565,0,Newman,0,0,Fiber Optic,37.343846,-121.039391,1,45.55,0,3,Offer B,8504,0,0,1,0,46,1,619.0,0.0,0.0,2062.15,0,0,95360
4522,1,0,1,0,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.7,587.1,0,45,0,22.89,2492,0,Oakdale,0,1,NA,37.785033,-120.776141,1,20.7,0,2,None,25384,0,0,1,0,30,0,0.0,686.7,0.0,587.1,0,0,95361
4523,1,1,1,0,10,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,75.3,720.45,0,80,30,25.13,4254,0,Patterson,0,1,DSL,37.410236,-121.32033700000001,1,75.3,0,7,None,15536,0,1,1,0,10,1,216.0,251.3,0.0,720.45,0,0,95363
4524,1,0,1,0,23,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,99.25,2186.4,1,33,8,19.2,5338,1,Pinecrest,1,1,Cable,38.224869,-119.755729,1,103.22,0,1,Offer D,235,0,1,1,0,23,2,175.0,441.6,0.0,2186.4,0,0,95364
4525,1,0,0,0,32,1,0,Fiber optic,1,1,0,1,Month-to-month,1,Credit card (automatic),93.4,2979.3,0,22,85,46.33,3224,0,Planada,1,1,Cable,37.329725,-120.306399,0,93.4,0,0,None,4150,0,0,0,1,32,1,2532.0,1482.56,0.0,2979.3,1,0,95365
4526,1,0,0,0,13,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),73.75,956.65,0,34,5,30.06,2070,0,Ripon,0,1,Fiber Optic,37.750778000000004,-121.13238,0,73.75,0,0,None,12646,0,0,0,0,13,1,4.78,390.78,0.0,956.65,0,1,95366
4527,0,0,0,0,39,1,0,Fiber optic,0,0,0,0,Two year,1,Electronic check,80.45,3201.55,1,39,30,24.45,2224,1,Riverbank,1,0,Fiber Optic,37.734971,-120.95427099999999,0,83.66799999999999,0,0,None,16525,1,1,0,0,39,2,960.0,953.55,0.0,3201.55,0,0,95367
4528,0,0,0,0,44,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),88.15,3973.2,0,35,24,32.83,4112,0,Salida,1,0,DSL,37.713152,-121.08738999999998,0,88.15,0,0,Offer B,12466,0,1,0,0,44,2,954.0,1444.52,0.0,3973.2,0,0,95368
4529,1,1,0,0,9,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,49.2,447.9,0,74,12,7.11,2145,0,Snelling,0,1,Fiber Optic,37.521708000000004,-120.42684299999999,0,49.2,0,0,None,1158,1,0,0,0,9,0,5.37,63.99,0.0,447.9,0,1,95369
4530,0,0,1,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.65,1335.2,0,22,0,33.01,4994,0,Sonora,0,0,NA,37.982715999999996,-120.343732,1,19.65,0,4,None,25340,0,0,1,0,67,1,0.0,2211.67,0.0,1335.2,1,0,95370
4531,1,0,1,1,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),79.35,661.25,1,30,65,31.67,4533,1,Soulsbyville,1,1,Cable,37.990574,-120.261821,1,82.524,0,1,None,1519,0,1,1,0,9,2,0.0,285.0300000000001,0.0,661.25,0,1,95372
4532,0,0,0,0,15,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.75,1111.85,1,42,23,42.83,2813,1,Stevinson,0,0,DSL,37.316807,-120.855753,0,82.94,0,0,Offer D,1960,0,0,0,0,15,1,256.0,642.4499999999998,0.0,1111.85,0,0,95374
4533,0,0,1,0,71,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),105.15,7555,0,37,3,10.46,5707,0,Tracy,1,0,Cable,37.680968,-121.446049,1,105.15,0,4,None,69801,0,0,1,1,71,0,0.0,742.6600000000002,0.0,7555.0,0,1,95376
4534,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),49.0,49,0,32,17,49.19,5289,0,Tuolumne,0,1,DSL,37.939768,-120.188002,0,49.0,0,0,None,3979,1,0,0,0,1,1,0.0,49.19,0.0,49.0,0,0,95379
4535,0,0,1,1,30,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.05,3046.15,1,64,24,39.74,4664,1,Turlock,1,0,DSL,37.474396,-120.87591699999999,1,104.052,0,1,None,40545,0,2,1,1,30,2,731.0,1192.2,0.0,3046.15,0,0,95380
4536,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.35,69.35,1,64,30,45.86,5796,1,Turlock,0,1,Fiber Optic,37.529656,-120.85435700000001,0,72.124,0,0,None,24708,0,0,0,0,1,1,0.0,45.86,0.0,69.35,0,1,95382
4537,1,0,1,0,17,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Mailed check,49.8,836.35,0,27,52,0.0,5575,0,Twain Harte,0,1,Fiber Optic,38.107440999999994,-120.230625,1,49.8,0,1,None,4848,0,0,1,1,17,1,0.0,0.0,0.0,836.35,1,1,95383
4538,0,0,0,0,3,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,85.8,272.2,1,20,80,10.6,5641,1,Vernalis,0,0,Fiber Optic,37.609095,-121.26338100000001,0,89.23200000000001,0,0,None,274,1,2,0,1,3,2,0.0,31.8,0.0,272.2,1,1,95385
4539,1,0,1,1,67,1,1,DSL,1,0,1,1,Two year,1,Electronic check,79.7,5293.4,1,49,3,42.77,6289,1,Waterford,1,1,DSL,37.669515999999994,-120.62696399999999,1,82.88799999999999,0,0,None,8308,0,0,0,1,67,2,0.0,2865.59,0.0,5293.4,0,1,95386
4540,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.95,20.95,0,52,0,2.29,2285,0,Escondido,0,1,NA,33.141265000000004,-116.967221,0,20.95,0,0,Offer E,48690,0,0,0,0,1,0,0.0,2.29,0.0,20.95,0,0,92027
4541,0,1,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.55,50.55,1,69,2,22.56,3357,1,Winton,0,0,Cable,37.421299,-120.59958700000001,0,52.572,0,0,None,11463,0,2,0,0,1,1,0.0,22.56,0.0,50.55,0,0,95388
4542,0,1,1,0,32,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,79.3,2570,0,68,11,2.17,5242,0,Escondido,1,0,Cable,33.141265000000004,-116.967221,1,79.3,0,2,Offer C,48690,0,0,1,0,32,1,283.0,69.44,0.0,2570.0,0,0,92027
4543,1,0,1,1,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.5,798.2,0,27,0,39.53,2446,0,Santa Rosa,0,1,NA,38.460516999999996,-122.79033500000001,1,19.5,1,8,Offer B,36125,0,0,1,0,41,1,0.0,1620.73,0.0,798.2,1,0,95401
4544,1,0,1,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.55,80.55,1,25,80,43.67,4273,1,Santa Rosa,0,1,Fiber Optic,38.488431,-122.752839,1,83.772,0,1,None,40270,0,1,1,1,1,2,0.0,43.67,0.0,80.55,1,1,95403
4545,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),44.15,44.15,0,45,13,9.82,3103,0,Santa Rosa,0,0,DSL,38.526941,-122.709096,0,44.15,0,0,Offer E,35057,0,0,0,0,1,0,0.0,9.82,0.0,44.15,0,0,95404
4546,0,0,1,1,12,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,84.5,916.9,1,28,65,40.63,4154,1,Santa Rosa,1,0,Cable,38.439696000000005,-122.66881699999999,1,87.88000000000002,0,1,None,22250,0,1,1,1,12,8,0.0,487.56000000000006,0.0,916.9,1,1,95405
4547,1,0,1,1,62,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,105.5,6487.2,0,22,52,14.75,4271,0,Santa Rosa,0,1,Fiber Optic,38.394090999999996,-122.739814,1,105.5,1,8,Offer B,30876,0,0,1,1,62,0,3373.0,914.5,0.0,6487.2,1,0,95407
4548,0,0,0,0,22,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Mailed check,84.3,1855.65,1,25,57,29.07,5313,1,Santa Rosa,0,0,Fiber Optic,38.468893,-122.58053899999999,0,87.67200000000001,0,0,None,25718,0,3,0,1,22,2,0.0,639.54,0.0,1855.65,1,1,95409
4549,0,0,0,1,17,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),92.7,1556.85,0,37,19,49.78,2347,0,Albion,1,0,Fiber Optic,39.225694,-123.717354,0,92.7,2,0,None,1054,1,0,0,0,17,2,0.0,846.26,0.0,1556.85,0,1,95410
4550,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),26.25,1988.05,0,37,0,2.57,5098,0,Annapolis,0,0,NA,38.731055,-123.316553,1,26.25,1,8,None,747,0,0,1,0,72,0,0.0,185.04,0.0,1988.05,0,0,95412
4551,1,0,1,1,56,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),96.95,5432.2,0,39,53,23.52,6484,0,Boonville,0,1,Cable,39.025867,-123.38154399999999,1,96.95,3,4,Offer B,1374,1,0,1,0,56,1,2879.0,1317.12,0.0,5432.2,0,0,95415
4552,0,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.45,147.55,0,32,0,45.99,2392,0,Branscomb,0,0,NA,39.710591,-123.682799,0,20.45,0,0,Offer E,176,0,0,0,0,9,0,0.0,413.91,0.0,147.55,0,0,95417
4553,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),115.8,8424.9,0,58,6,43.12,6479,0,Caspar,1,1,Fiber Optic,39.361283,-123.784599,1,115.8,0,0,None,333,1,0,0,1,72,0,505.0,3104.64,0.0,8424.9,0,0,95420
4554,1,0,0,0,20,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),108.2,2203.7,0,40,18,16.05,2102,0,Cazadero,1,1,Fiber Optic,38.578807,-123.19338,0,108.2,0,0,None,1575,1,0,0,1,20,0,397.0,321.0,0.0,2203.7,0,0,95421
4555,1,0,1,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.2,387.4,0,32,0,31.7,4821,0,Clearlake,0,1,NA,38.965804,-122.63177900000001,1,20.2,3,3,None,13485,0,0,1,0,19,0,0.0,602.3,0.0,387.4,0,0,95422
4556,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,67.75,116.65,1,58,4,11.75,2299,1,Clearlake Oaks,0,1,Fiber Optic,39.07116,-122.598542,0,70.46000000000002,0,0,None,3684,0,0,0,0,2,2,5.0,23.5,0.0,116.65,0,0,95423
4557,1,0,0,0,53,0,No phone service,DSL,0,0,1,1,One year,0,Credit card (automatic),54.9,3045.75,0,62,17,0.0,5677,0,Cloverdale,1,1,Fiber Optic,38.801936,-122.93893500000001,0,54.9,0,0,Offer B,9210,1,0,0,1,53,2,0.0,0.0,0.0,3045.75,0,1,95425
4558,0,1,0,0,27,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.25,2287.25,1,74,28,31.17,5172,1,Cobb,0,0,Fiber Optic,38.838088,-122.73203000000001,0,88.66,0,0,None,1591,0,2,0,1,27,7,640.0,841.59,0.0,2287.25,0,0,95426
4559,1,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.15,130.5,0,56,0,6.93,5761,0,Comptche,0,1,NA,39.239818,-123.565432,0,20.15,0,0,None,371,0,0,0,0,6,2,0.0,41.58,0.0,130.5,0,0,95427
4560,1,0,1,1,9,1,1,Fiber optic,0,0,1,0,One year,1,Electronic check,90.35,767.9,0,22,82,30.46,2993,0,Covelo,1,1,Fiber Optic,39.83307,-123.17876499999998,1,90.35,3,9,Offer E,2296,0,0,1,0,9,2,630.0,274.14,0.0,767.9,1,0,95428
4561,0,0,1,1,8,1,1,DSL,0,1,0,0,Month-to-month,0,Electronic check,55.75,446.8,0,62,53,12.41,5681,0,Dos Rios,0,0,Cable,39.756049,-123.358701,1,55.75,3,1,Offer E,91,0,0,1,0,8,0,0.0,99.28,0.0,446.8,0,1,95429
4562,0,0,1,1,71,1,1,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),114.6,8100.25,0,45,29,4.91,4071,0,Duncans Mills,1,0,Fiber Optic,38.445603000000006,-123.06375600000001,1,114.6,3,5,None,187,1,0,1,1,71,2,0.0,348.61,0.0,8100.25,0,1,95430
4563,0,0,0,0,10,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.05,830.7,1,60,11,49.7,3740,1,Eldridge,0,0,DSL,38.348884000000005,-122.51698999999999,0,83.25200000000001,0,0,None,363,0,0,0,0,10,3,91.0,497.0,0.0,830.7,0,0,95431
4564,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,20,1,30,0,46.77,3657,1,Elk,0,1,NA,39.108252,-123.645121,0,20.0,0,0,None,383,0,0,0,0,1,3,0.0,46.77,0.0,20.0,0,0,95432
4565,0,0,1,0,71,0,No phone service,DSL,1,1,1,1,One year,0,Bank transfer (automatic),66.8,4689.15,0,23,85,0.0,4698,0,Forestville,1,0,DSL,38.499302,-122.92443999999999,1,66.8,0,10,None,6216,1,0,1,1,71,1,3986.0,0.0,0.0,4689.15,1,0,95436
4566,1,0,1,0,68,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,100.3,6754.35,0,43,3,49.51,5757,0,Fort Bragg,0,1,Fiber Optic,39.455555,-123.68397900000001,1,100.3,0,1,None,14417,1,0,1,1,68,2,203.0,3366.68,0.0,6754.35,0,0,95437
4567,1,0,0,0,34,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.35,3540.65,0,51,18,28.0,5503,0,Fulton,0,1,Cable,38.493888,-122.77714099999999,0,105.35,0,0,None,476,1,0,0,1,34,0,0.0,952.0,0.0,3540.65,0,1,95439
4568,1,0,0,0,26,1,0,Fiber optic,0,1,0,0,One year,1,Electronic check,85.2,2184.6,0,51,11,29.72,5156,0,Geyserville,1,1,Fiber Optic,38.731771,-123.064272,0,85.2,0,0,None,2349,1,0,0,0,26,2,240.0,772.72,0.0,2184.6,0,0,95441
4569,0,0,0,0,22,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),48.8,1054.6,1,32,33,3.95,2270,1,Glen Ellen,0,0,Cable,38.368744,-122.52264199999999,0,50.752,0,0,None,4101,0,0,0,0,22,0,34.8,86.9,0.0,1054.6,0,1,95442
4570,1,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,18.95,130.55,0,42,0,33.18,4097,0,Glenhaven,0,1,NA,39.045246,-122.743181,0,18.95,0,0,Offer E,175,0,0,0,0,7,1,0.0,232.26,0.0,130.55,0,0,95443
4571,0,0,1,0,20,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.8,1540.35,0,51,28,43.49,5456,0,Graton,0,0,Fiber Optic,38.434362,-122.86891000000001,1,69.8,0,0,None,390,0,0,0,0,20,2,0.0,869.8000000000002,0.0,1540.35,0,1,95444
4572,0,0,1,0,60,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.15,6411.25,0,48,22,9.98,4115,0,Gualala,1,0,Fiber Optic,38.848082,-123.50608000000001,1,106.15,0,5,Offer B,1916,0,0,1,1,60,1,0.0,598.8000000000002,0.0,6411.25,0,1,95445
4573,1,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,20.55,1432.55,0,51,0,37.11,5809,0,Guerneville,0,1,NA,38.52576,-123.013347,1,20.55,1,5,None,4913,0,0,1,0,72,1,0.0,2671.92,0.0,1432.55,0,0,95446
4574,0,1,1,0,72,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),105.75,7629.85,0,70,16,18.15,5832,0,Healdsburg,1,0,Fiber Optic,38.618347,-122.908422,1,105.75,0,7,Offer A,17979,0,0,1,1,72,0,0.0,1306.8,0.0,7629.85,0,1,95448
4575,1,0,0,0,4,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,25.25,101.9,0,64,0,3.69,3962,0,Hopland,0,1,NA,38.937059999999995,-123.11811100000001,0,25.25,0,0,Offer E,1373,0,1,0,0,4,2,0.0,14.76,0.0,101.9,0,0,95449
4576,1,0,1,1,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.75,313.4,0,40,0,31.99,3677,0,Jenner,0,1,NA,38.505995,-123.18701899999999,1,19.75,1,2,None,438,0,0,1,0,16,0,0.0,511.84,0.0,313.4,0,0,95450
4577,0,1,1,0,62,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,104.85,6312.9,0,70,18,22.74,5061,0,Kelseyville,1,0,Cable,38.93496,-122.792243,1,104.85,0,8,Offer B,9902,0,0,1,1,62,2,0.0,1409.88,0.0,6312.9,0,1,95451
4578,0,0,0,0,10,1,0,DSL,0,0,0,1,Month-to-month,1,Mailed check,60.95,629.55,0,58,29,8.35,4323,0,Kenwood,0,0,DSL,38.419525,-122.52158500000002,0,60.95,0,0,None,1653,1,0,0,1,10,0,0.0,83.5,0.0,629.55,0,1,95452
4579,1,0,0,0,31,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,81.15,2640.55,0,60,12,42.05,3031,0,Lakeport,0,1,Cable,39.080469,-122.955176,0,81.15,0,0,None,11180,0,0,0,0,31,0,0.0,1303.55,0.0,2640.55,0,1,95453
4580,0,0,1,0,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.1,1372.45,0,26,0,39.44,4241,0,Laytonville,0,0,NA,39.806141,-123.531098,1,19.1,0,2,None,2706,0,0,1,0,71,0,0.0,2800.24,0.0,1372.45,1,0,95454
4581,1,0,0,0,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.8,1212.25,0,29,0,49.02,4758,0,Little River,0,1,NA,39.245911,-123.77214,0,20.8,0,0,Offer B,882,0,1,0,0,58,1,0.0,2843.1600000000008,0.0,1212.25,1,0,95456
4582,1,0,1,1,70,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),90.15,6237.05,0,31,13,2.5,5824,0,Lower Lake,1,1,Fiber Optic,38.925545,-122.54908300000001,1,90.15,1,7,None,2644,1,0,1,1,70,0,81.08,175.0,0.0,6237.05,0,1,95457
4583,0,0,1,0,71,1,1,DSL,1,1,1,1,Two year,0,Electronic check,90.1,6310.9,0,30,71,22.33,5054,0,Lucerne,1,0,DSL,39.141934,-122.770679,1,90.1,0,2,None,3002,1,0,1,1,71,1,4481.0,1585.4299999999996,0.0,6310.9,0,0,95458
4584,1,1,0,0,69,1,1,DSL,1,0,0,1,Two year,0,Credit card (automatic),74.1,5031,0,71,10,13.36,4204,0,Manchester,1,1,Cable,38.966713,-123.58641200000001,0,74.1,0,0,Offer A,586,1,0,0,1,69,0,503.0,921.84,0.0,5031.0,0,0,95459
4585,0,1,0,0,1,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.05,85.05,1,68,8,16.37,2975,1,Mendocino,0,0,Cable,39.305545,-123.743697,0,88.45200000000001,0,0,None,2229,0,1,0,1,1,3,0.0,16.37,0.0,85.05,0,0,95460
4586,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),118.75,8672.45,0,33,53,41.14,5475,0,Middletown,1,0,DSL,38.787446,-122.58675,1,118.75,3,1,None,7789,1,0,1,1,72,1,0.0,2962.08,0.0,8672.45,0,1,95461
4587,0,0,1,0,26,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Credit card (automatic),85.9,2196.45,0,56,2,42.26,4038,0,Monte Rio,0,0,Cable,38.471049,-123.015549,1,85.9,0,1,None,1537,1,0,1,1,26,0,0.0,1098.76,0.0,2196.45,0,1,95462
4588,0,0,1,0,33,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),95.0,3008.15,0,41,22,10.34,4639,0,Navarro,1,0,DSL,39.182916,-123.552571,1,95.0,0,1,None,148,1,0,1,1,33,0,0.0,341.22,0.0,3008.15,0,1,95463
4589,0,0,1,1,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.15,220.8,0,51,0,18.62,2836,0,Nice,0,0,NA,39.12334,-122.83819799999999,1,20.15,3,1,None,2223,0,0,1,0,10,1,0.0,186.2,0.0,220.8,0,0,95464
4590,0,1,0,0,57,1,1,Fiber optic,1,0,0,1,Two year,0,Credit card (automatic),101.3,5779.6,0,80,17,36.89,4421,0,Occidental,1,0,DSL,38.415003000000006,-122.998726,0,101.3,0,0,Offer B,1880,1,0,0,1,57,1,983.0,2102.73,0.0,5779.6,0,0,95465
4591,0,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,21.2,222.65,0,52,0,10.46,2066,0,Philo,0,0,NA,39.094102,-123.500853,0,21.2,0,0,None,1113,0,0,0,0,10,0,0.0,104.6,0.0,222.65,0,0,95466
4592,0,0,1,1,39,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,24.2,914.6,0,31,0,5.88,3109,0,Point Arena,0,0,NA,38.911299,-123.60958799999999,1,24.2,2,1,None,1352,0,0,1,0,39,2,0.0,229.32,0.0,914.6,0,0,95468
4593,0,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.3,246.3,0,40,0,48.92,4188,0,Potter Valley,0,0,NA,39.408634,-123.04551599999999,0,20.3,0,0,None,1884,0,0,0,0,11,1,0.0,538.12,0.0,246.3,0,0,95469
4594,0,0,1,1,21,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,102.8,2110.15,1,52,3,16.67,3123,1,Redwood Valley,1,0,Fiber Optic,39.298065,-123.25211000000002,1,106.912,0,1,None,5995,1,3,1,1,21,1,63.0,350.07000000000005,0.0,2110.15,0,0,95470
4595,0,0,1,1,68,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),85.3,5560,0,36,26,25.16,4732,0,Rio Nido,1,0,Fiber Optic,38.522328,-122.97932,1,85.3,2,1,None,298,1,0,1,1,68,1,1446.0,1710.88,0.0,5560.0,0,0,95471
4596,1,0,0,0,18,1,1,Fiber optic,0,0,1,0,One year,1,Credit card (automatic),89.6,1633,0,43,2,34.78,2269,0,Sebastopol,1,1,Fiber Optic,38.398815,-122.861923,0,89.6,0,0,None,31266,0,0,0,0,18,0,0.0,626.04,0.0,1633.0,0,1,95472
4597,0,0,0,0,6,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,99.95,547.65,1,26,65,5.16,3722,1,Sonoma,1,0,DSL,38.25485,-122.461799,0,103.948,0,0,None,34314,1,1,0,1,6,3,0.0,30.96,0.0,547.65,1,1,95476
4598,1,0,0,0,18,1,1,DSL,1,0,0,0,Month-to-month,0,Mailed check,56.25,969.85,0,47,17,33.8,2277,0,Ukiah,0,1,Fiber Optic,39.134075,-123.23422,0,56.25,0,0,None,30988,0,0,0,0,18,0,0.0,608.4,0.0,969.85,0,1,95482
4599,0,0,1,1,52,1,0,DSL,0,0,0,0,One year,1,Bank transfer (automatic),50.95,2610.65,0,59,29,10.03,4298,0,Upper Lake,1,0,Fiber Optic,39.220368,-122.907693,1,50.95,2,2,Offer B,2344,0,0,1,0,52,1,0.0,521.56,0.0,2610.65,0,1,95485
4600,1,0,1,1,56,1,1,Fiber optic,1,1,1,1,Two year,0,Mailed check,115.85,6567.9,0,42,27,40.86,4937,0,Westport,1,1,Fiber Optic,39.724433000000005,-123.767578,1,115.85,3,8,Offer B,309,1,1,1,1,56,1,0.0,2288.16,0.0,6567.9,0,1,95488
4601,1,0,0,0,45,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),103.65,4747.85,0,51,13,24.75,2183,0,Willits,1,1,DSL,39.492046,-123.375818,0,103.65,0,0,Offer B,13472,1,0,0,1,45,2,0.0,1113.75,0.0,4747.85,0,1,95490
4602,0,0,0,0,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,26.1,1759.55,0,45,0,43.3,6466,0,Windsor,0,0,NA,38.527297,-122.81004399999999,0,26.1,0,0,None,23701,0,0,0,0,67,0,0.0,2901.1,0.0,1759.55,0,0,95492
4603,1,0,1,0,3,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,35.1,101.1,0,33,25,0.0,3610,0,Witter Springs,0,1,Fiber Optic,39.222322999999996,-122.98548799999999,1,35.1,0,3,Offer E,240,1,0,1,0,3,2,0.0,0.0,0.0,101.1,0,1,95493
4604,1,1,0,0,65,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),99.1,6496.15,0,80,3,18.23,4574,0,Yorkville,1,1,DSL,38.888351,-123.23964699999999,0,99.1,0,0,Offer B,335,0,0,0,1,65,2,0.0,1184.95,0.0,6496.15,0,1,95494
4605,1,0,1,0,63,1,1,DSL,0,1,0,1,Two year,0,Mailed check,67.25,4234.15,0,52,28,48.14,6438,0,The Sea Ranch,0,1,Cable,38.696659000000004,-123.43686100000001,1,67.25,0,2,None,752,1,0,1,1,63,2,1186.0,3032.82,0.0,4234.15,0,0,95497
4606,0,0,1,1,11,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.0,300.7,0,50,0,15.04,5409,0,Eureka,0,0,NA,40.796621,-124.15428,1,25.0,2,1,None,23224,0,0,1,0,11,2,0.0,165.44,0.0,300.7,0,0,95501
4607,1,0,0,1,1,1,0,DSL,0,0,0,1,Month-to-month,1,Mailed check,59.55,59.55,0,20,48,41.39,5824,0,Eureka,0,1,Fiber Optic,40.737431,-124.108897,0,59.55,1,0,None,23570,1,0,0,1,1,0,0.0,41.39,0.0,59.55,1,0,95503
4608,1,0,0,0,55,1,1,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),77.8,4323.35,0,48,23,26.3,6483,0,Alderpoint,1,1,Fiber Optic,40.166028000000004,-123.584144,0,77.8,0,0,None,261,0,0,0,1,55,0,994.0,1446.5,0.0,4323.35,0,0,95511
4609,1,0,1,1,25,1,1,DSL,0,0,0,0,One year,1,Mailed check,55.1,1466.1,0,34,25,47.1,2499,0,Blocksburg,0,1,Cable,40.309088,-123.668201,1,55.1,1,2,None,199,1,0,1,0,25,1,0.0,1177.5,0.0,1466.1,0,1,95514
4610,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),117.8,8684.8,1,31,9,34.87,4432,1,Mckinleyville,1,1,Fiber Optic,40.965011,-124.01525500000001,1,122.512,0,1,None,15921,1,1,1,1,72,1,0.0,2510.64,0.0,8684.8,0,1,95519
4611,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.15,1776.45,0,55,0,37.98,5613,0,Arcata,0,0,NA,40.839958,-124.00375700000001,1,24.15,0,7,None,19596,0,0,1,0,72,0,0.0,2734.56,0.0,1776.45,0,0,95521
4612,0,0,0,1,65,0,No phone service,DSL,0,1,1,0,Two year,0,Mailed check,45.25,2933.95,0,33,25,0.0,5712,0,Bayside,0,0,Fiber Optic,40.825486,-124.049485,0,45.25,2,0,None,1689,1,0,0,0,65,0,73.35,0.0,0.0,2933.95,0,1,95524
4613,0,1,0,0,54,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.5,4370.25,1,68,11,45.77,5684,1,Blue Lake,0,0,DSL,40.94338,-123.831799,0,82.68,0,0,None,1584,0,1,0,0,54,5,481.0,2471.580000000001,0.0,4370.25,0,0,95525
4614,1,0,1,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,144.35,0,31,0,39.98,4954,0,Bridgeville,0,1,NA,40.372532,-123.525626,1,20.25,1,9,None,695,0,0,1,0,7,1,0.0,279.86,0.0,144.35,0,0,95526
4615,0,0,1,0,72,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),64.75,4804.75,0,45,26,15.23,4675,0,Burnt Ranch,0,0,Cable,40.854512,-123.450097,1,64.75,0,7,None,485,1,0,1,0,72,1,1249.0,1096.56,0.0,4804.75,0,0,95527
4616,1,0,1,0,21,1,0,DSL,0,0,1,0,Month-to-month,0,Bank transfer (automatic),54.6,1125.2,0,57,11,17.19,5763,0,Carlotta,0,1,Fiber Optic,40.497283,-123.93037,1,54.6,0,4,None,1072,0,0,1,0,21,0,124.0,360.99,0.0,1125.2,0,0,95528
4617,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.7,39.85,0,28,0,13.89,2107,0,Fallbrook,0,0,NA,33.362575,-117.299644,0,20.7,0,0,None,42239,0,0,0,0,2,0,0.0,27.78,0.0,39.85,1,0,92028
4618,1,1,0,0,4,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.75,422.4,0,80,17,19.0,2757,0,Ferndale,1,1,DSL,40.4785,-124.301372,0,94.75,0,0,None,2965,0,0,0,1,4,0,0.0,76.0,0.0,422.4,0,1,95536
4619,1,0,1,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),79.65,251.75,1,33,19,43.27,5036,1,Fields Landing,0,1,Cable,40.726949,-124.217378,1,82.83600000000001,0,1,None,228,1,0,1,0,3,0,48.0,129.81,0.0,251.75,0,0,95537
4620,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),115.8,8332.15,0,50,25,27.59,5130,0,Fortuna,1,1,DSL,40.584990999999995,-124.121504,1,115.8,0,8,None,12241,1,0,1,1,72,1,0.0,1986.48,0.0,8332.15,0,1,95540
4621,0,0,0,0,6,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.45,314.6,0,63,8,39.16,3672,0,Garberville,0,0,Fiber Optic,40.057784000000005,-123.679461,0,49.45,0,0,None,2423,0,0,0,0,6,1,0.0,234.96,0.0,314.6,0,1,95542
4622,1,0,0,0,52,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),83.8,4331.4,0,58,23,5.92,6339,0,Gasquet,1,1,Cable,41.867908,-123.79414399999999,0,83.8,0,0,None,532,0,0,0,1,52,0,996.0,307.84,0.0,4331.4,0,0,95543
4623,1,1,1,0,69,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),95.35,6382,0,73,13,49.91,6132,0,Honeydew,1,1,Fiber Optic,40.342928,-124.06332900000001,1,95.35,0,5,None,82,0,0,1,1,69,3,830.0,3443.79,0.0,6382.0,0,0,95545
4624,1,0,0,0,8,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.7,740.3,1,44,11,19.49,5811,1,Hoopa,1,1,DSL,41.163637,-123.70484099999999,0,98.488,0,0,None,3041,0,0,0,1,8,0,81.0,155.92,0.0,740.3,0,0,95546
4625,0,1,0,0,8,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.05,600.15,0,72,13,2.18,4899,0,Hydesville,1,0,Fiber Optic,40.557314,-124.08166200000001,0,74.05,0,0,None,1201,0,0,0,0,8,1,0.0,17.44,0.0,600.15,0,1,95547
4626,0,1,0,0,63,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),89.6,5538.8,0,74,16,41.8,4438,0,Klamath,1,0,DSL,41.572813000000004,-124.03501100000001,0,89.6,0,0,Offer B,1215,0,0,0,1,63,0,0.0,2633.4,0.0,5538.8,0,1,95548
4627,1,0,0,0,60,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),116.6,7049.5,0,22,52,44.24,5680,0,Kneeland,1,1,Cable,40.664483000000004,-123.865325,0,116.6,0,0,None,264,1,0,0,1,60,2,3666.0,2654.4,0.0,7049.5,1,0,95549
4628,0,0,1,0,12,1,0,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),54.2,690.5,0,24,51,23.99,4474,0,Korbel,0,0,Fiber Optic,40.7666,-123.80458,1,54.2,0,4,Offer D,155,1,0,1,0,12,1,0.0,287.88,0.0,690.5,1,1,95550
4629,0,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.3,279.3,0,50,0,21.36,5917,0,Loleta,0,0,NA,40.665952000000004,-124.240051,0,19.3,0,0,Offer D,1447,0,0,0,0,13,1,0.0,277.68,0.0,279.3,0,0,95551
4630,1,0,0,0,22,1,1,DSL,1,1,0,0,Month-to-month,0,Mailed check,65.05,1427.55,0,20,47,43.78,4709,0,Mad River,1,1,Fiber Optic,40.390301,-123.412327,0,65.05,0,0,Offer D,265,0,0,0,0,22,1,0.0,963.16,0.0,1427.55,1,1,95552
4631,1,0,0,0,5,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,92.5,452.7,1,33,28,3.25,2810,1,Miranda,1,1,Cable,40.210895,-123.86,0,96.2,0,0,None,867,0,0,0,0,5,0,127.0,16.25,0.0,452.7,0,0,95553
4632,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.45,19.45,1,54,0,28.73,2865,1,Myers Flat,0,0,NA,40.267158,-123.80591299999999,1,19.45,2,1,None,644,0,2,1,0,1,1,0.0,28.73,0.0,19.45,0,0,95554
4633,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.05,1709.15,0,59,0,48.29,4755,0,Orick,0,0,NA,41.336354,-124.044354,1,24.05,3,4,None,494,0,0,1,0,72,2,0.0,3476.88,0.0,1709.15,0,0,95555
4634,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),18.75,53.15,0,23,0,4.92,5355,0,Orleans,0,0,NA,41.269521000000005,-123.546958,0,18.75,0,0,None,574,0,1,0,0,2,3,0.0,9.84,0.0,53.15,1,0,95556
4635,0,0,1,1,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.15,777.35,0,42,0,3.01,3556,0,Petrolia,0,0,NA,40.274302,-124.210902,1,20.15,3,1,None,300,0,1,1,0,40,1,0.0,120.4,0.0,777.35,0,0,95558
4636,1,0,1,1,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.0,860.85,0,23,0,36.86,3743,0,Phillipsville,0,1,NA,40.184094,-123.74548700000001,1,20.0,3,2,None,163,0,0,1,0,44,0,0.0,1621.84,0.0,860.85,1,0,95559
4637,1,1,1,0,71,1,0,DSL,1,1,1,0,One year,1,Bank transfer (automatic),71.0,5012.1,0,69,24,11.35,5247,0,Redway,0,1,DSL,40.142256,-123.85292700000001,1,71.0,0,10,None,1851,1,0,1,0,71,0,0.0,805.85,0.0,5012.1,0,1,95560
4638,0,0,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.55,166.3,1,32,31,41.37,4320,1,Rio Dell,0,0,Fiber Optic,40.485849,-124.163234,0,78.572,0,0,None,3284,0,0,0,0,2,1,52.0,82.74,0.0,166.3,0,0,95562
4639,1,1,0,0,26,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.6,2404.1,0,65,9,25.04,4030,0,Salyer,0,1,DSL,40.89866,-123.539754,0,93.6,0,0,Offer C,660,0,0,0,1,26,1,216.0,651.04,0.0,2404.1,0,0,95563
4640,1,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.0,70,1,38,4,38.8,2485,1,Samoa,0,1,DSL,40.809636,-124.189977,1,72.8,0,1,None,395,0,1,1,0,1,2,0.0,38.8,0.0,70.0,0,0,95564
4641,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,24.4,24.4,0,19,76,0.0,5092,0,Scotia,0,0,DSL,40.440636,-124.098739,0,24.4,0,0,None,1125,0,0,0,1,1,0,0.0,0.0,0.0,24.4,1,1,95565
4642,1,0,1,1,65,1,0,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),74.8,4820.15,1,56,33,40.47,5207,1,Smith River,0,1,DSL,41.950683000000005,-124.097094,1,77.792,0,1,Offer B,2020,1,3,1,1,65,5,1591.0,2630.55,0.0,4820.15,0,0,95567
4643,1,0,0,0,3,1,1,DSL,0,0,1,0,Month-to-month,1,Mailed check,65.25,209.9,0,32,27,42.68,2562,0,Somes Bar,0,1,Fiber Optic,41.444606,-123.47189499999999,0,65.25,0,0,None,202,1,2,0,0,3,2,0.0,128.04,0.0,209.9,0,1,95568
4644,1,0,0,0,13,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.55,610.75,0,28,59,33.95,5530,0,Redcrest,0,1,Fiber Optic,40.363446,-123.83504099999999,0,50.55,0,0,Offer D,400,1,0,0,1,13,0,0.0,441.35,0.0,610.75,1,1,95569
4645,0,0,1,0,33,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.4,3409.6,1,46,13,11.32,3185,1,Trinidad,1,0,DSL,41.162295,-124.027381,1,108.576,0,1,None,2369,0,3,1,1,33,2,443.0,373.56,0.0,3409.6,0,0,95570
4646,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.7,70.7,0,19,52,38.81,4056,0,Weott,0,0,DSL,40.310119,-123.909449,0,70.7,0,0,None,270,0,0,0,1,1,3,0.0,38.81,0.0,70.7,1,0,95571
4647,1,0,1,1,4,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.25,155.35,0,33,30,35.09,2776,0,Willow Creek,0,1,DSL,40.949011999999996,-123.655847,1,45.25,2,8,Offer E,1666,0,0,1,0,4,1,47.0,140.36,0.0,155.35,0,0,95573
4648,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,144,0,51,26,1.57,2980,0,Leggett,0,1,DSL,39.873371,-123.741474,0,70.3,0,0,Offer E,321,0,0,0,0,2,1,0.0,3.14,0.0,144.0,0,1,95585
4649,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),108.95,7875,0,28,53,21.26,5758,0,Piercy,0,1,Cable,39.955587,-123.681175,1,108.95,0,0,None,200,1,0,0,1,72,1,0.0,1530.72,0.0,7875.0,1,1,95587
4650,0,0,1,1,37,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,26.45,911.6,0,42,0,31.83,5359,0,Fallbrook,0,0,NA,33.362575,-117.299644,1,26.45,2,1,None,42239,0,0,1,0,37,1,0.0,1177.71,0.0,911.6,0,0,92028
4651,0,0,0,0,15,1,0,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,86.2,1270.2,1,21,65,20.03,5829,1,Zenia,0,0,DSL,40.170357,-123.417298,0,89.64800000000002,0,0,None,259,0,0,0,1,15,4,826.0,300.4500000000001,0.0,1270.2,1,0,95595
4652,0,0,0,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),19.65,478.1,0,34,0,10.41,5916,0,Amador City,0,0,NA,38.431407,-120.8421,0,19.65,0,0,Offer D,222,0,0,0,0,23,0,0.0,239.43,0.0,478.1,0,0,95601
4653,0,0,1,1,30,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Credit card (automatic),51.2,1561.5,1,57,13,0.0,4568,1,Auburn,0,0,Cable,38.99003,-121.11440800000001,1,53.24800000000001,2,1,None,18197,1,1,1,1,30,6,203.0,0.0,0.0,1561.5,0,0,95602
4654,0,0,1,1,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,19.05,761.85,0,31,0,34.66,5091,0,Auburn,0,0,NA,38.912881,-121.08276599999999,1,19.05,3,4,None,24944,0,0,1,0,42,1,0.0,1455.7199999999998,0.0,761.85,0,0,95603
4655,0,0,0,0,32,1,1,DSL,1,0,1,1,One year,0,Mailed check,74.75,2282.95,0,45,5,33.45,2830,0,West Sacramento,0,0,Fiber Optic,38.592745,-121.54003600000001,0,74.75,0,0,Offer C,12756,0,0,0,1,32,1,0.0,1070.4,0.0,2282.95,0,1,95605
4656,0,0,1,1,22,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.8,1615.1,0,59,58,4.67,4479,0,Brooks,0,0,Fiber Optic,38.809804,-122.24138300000001,1,75.8,3,3,Offer D,382,0,0,1,0,22,0,937.0,102.74,0.0,1615.1,0,0,95606
4657,1,0,1,0,42,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),25.1,1097.15,0,26,59,0.0,4959,0,Capay,0,1,Fiber Optic,38.681651,-122.130569,1,25.1,0,5,None,262,0,0,1,1,42,2,647.0,0.0,0.0,1097.15,1,0,95607
4658,0,0,0,0,8,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.45,369.3,0,56,16,10.91,4909,0,Carmichael,0,0,Cable,38.626128,-121.328011,0,44.45,0,0,None,58830,0,0,0,0,8,0,5.91,87.28,0.0,369.3,0,1,95608
4659,0,0,1,1,65,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),104.3,6725.3,0,23,59,13.17,4997,0,Citrus Heights,1,0,Fiber Optic,38.69508,-121.271616,1,104.3,1,5,None,43718,0,0,1,1,65,1,3968.0,856.05,0.0,6725.3,1,0,95610
4660,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.5,31.55,1,23,0,28.02,2484,1,Clarksburg,0,0,NA,38.384648,-121.578701,0,19.5,0,0,None,1417,0,1,0,0,2,4,0.0,56.04,0.0,31.55,1,0,95612
4661,0,0,1,1,70,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),89.0,6293.2,0,30,51,33.24,5650,0,Cool,1,0,Cable,38.880621999999995,-120.97386499999999,1,89.0,1,3,None,3674,1,0,1,1,70,0,0.0,2326.8,0.0,6293.2,0,1,95614
4662,1,0,0,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.15,432.5,0,43,0,34.07,2722,0,Courtland,0,1,NA,38.311609000000004,-121.554034,0,20.15,2,0,Offer D,699,0,0,0,0,22,3,0.0,749.54,0.0,432.5,0,0,95615
4663,0,1,0,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.9,321.75,1,68,32,26.23,2122,1,Davis,0,0,Cable,38.508734999999994,-121.67881299999999,0,77.89600000000002,0,0,None,67411,0,0,0,0,4,2,103.0,104.92,0.0,321.75,0,0,95616
4664,0,0,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),74.9,147.15,1,37,20,38.28,2078,1,Davis,0,0,Fiber Optic,38.544002,-121.68555900000001,0,77.89600000000002,0,0,None,648,0,1,0,0,2,5,29.0,76.56,0.0,147.15,0,0,95618
4665,0,0,1,1,67,0,No phone service,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),36.15,2434.45,0,58,15,0.0,6314,0,Diamond Springs,0,0,DSL,38.683605,-120.811852,1,36.15,1,5,None,4426,0,0,1,0,67,0,365.0,0.0,0.0,2434.45,0,0,95619
4666,0,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.2,532.1,0,42,0,6.0,2159,0,Dixon,0,0,NA,38.392821000000005,-121.799917,0,19.2,0,0,Offer C,18529,0,0,0,0,25,2,0.0,150.0,0.0,532.1,0,0,95620
4667,0,0,1,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.25,375.25,0,49,0,48.03,4137,0,Citrus Heights,0,0,NA,38.69549,-121.307864,1,19.25,0,0,Offer D,41636,0,0,0,0,20,1,0.0,960.6,0.0,375.25,0,0,95621
4668,0,0,0,1,2,1,0,DSL,1,0,0,1,Month-to-month,1,Credit card (automatic),61.2,125.95,0,28,52,32.06,5056,0,El Dorado,0,0,DSL,38.63153,-120.84260900000001,0,61.2,2,0,Offer E,4097,0,0,0,1,2,2,0.0,64.12,0.0,125.95,1,1,95623
4669,1,0,0,0,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.45,1042.65,0,36,0,47.43,6097,0,Elk Grove,0,1,NA,38.434138,-121.30587,0,20.45,0,0,None,38534,0,0,0,0,51,0,0.0,2418.93,0.0,1042.65,0,0,95624
4670,0,0,1,1,46,0,No phone service,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),35.05,1620.25,0,27,52,0.0,4829,0,Elmira,0,0,Fiber Optic,38.349195,-121.902943,1,35.05,2,9,None,171,0,0,1,1,46,0,843.0,0.0,0.0,1620.25,1,0,95625
4671,0,0,0,0,25,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.25,2387.75,1,59,3,36.24,2195,1,Elverta,0,0,DSL,38.734997,-121.463719,0,104.26,0,0,None,6197,0,0,0,1,25,4,72.0,906.0,0.0,2387.75,0,0,95626
4672,1,0,0,1,13,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.0,659.35,0,20,27,26.63,5611,0,Esparto,0,1,Fiber Optic,38.834469,-122.12719299999999,0,44.0,1,0,Offer D,2756,0,0,0,1,13,0,0.0,346.19,0.0,659.35,1,1,95627
4673,0,1,0,0,25,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Mailed check,102.8,2660.2,1,75,33,36.5,4969,1,Fair Oaks,0,0,Cable,38.652065,-121.25441000000001,0,106.912,0,0,None,40750,0,0,0,0,25,3,878.0,912.5,0.0,2660.2,0,0,95628
4674,1,0,1,1,26,1,0,DSL,0,0,0,0,One year,0,Mailed check,50.35,1285.8,0,32,19,4.62,3386,0,Fiddletown,1,1,DSL,38.513484000000005,-120.704613,1,50.35,1,4,Offer C,850,0,0,1,0,26,1,0.0,120.12,0.0,1285.8,0,1,95629
4675,1,0,0,0,43,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,100.0,4211.55,1,56,25,39.37,4760,1,Folsom,0,1,DSL,38.672638,-121.147403,0,104.0,0,0,Offer B,51855,1,0,0,1,43,0,1053.0,1692.91,0.0,4211.55,0,0,95630
4676,1,0,0,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.0,377.55,0,41,0,24.1,5188,0,Foresthill,0,1,NA,39.031876000000004,-120.81114099999999,0,20.0,3,0,Offer D,5714,0,0,0,0,19,1,0.0,457.9,0.0,377.55,0,0,95631
4677,1,0,1,0,10,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.85,990.9,1,58,13,43.28,4243,1,Galt,0,1,DSL,38.274451,-121.259201,1,103.844,0,5,None,24194,1,4,1,1,10,1,0.0,432.8,0.0,990.9,0,1,95632
4678,0,0,0,1,2,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),94.2,193.8,1,34,14,42.89,5299,1,Garden Valley,0,0,DSL,38.852544,-120.83766899999999,0,97.96799999999999,0,0,None,2536,0,1,0,1,2,5,0.0,85.78,0.0,193.8,0,1,95633
4679,0,0,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),86.4,6058.95,0,21,41,15.35,6114,0,Georgetown,0,0,Fiber Optic,38.9386,-120.78551399999999,1,86.4,0,6,None,2723,1,0,1,1,72,0,248.42,1105.2,0.0,6058.95,1,1,95634
4680,1,1,0,0,18,1,1,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),58.4,964.9,0,73,7,47.34,2812,0,Greenwood,0,1,Fiber Optic,38.921333000000004,-120.897718,0,58.4,0,0,Offer D,1140,0,0,0,0,18,1,68.0,852.1200000000001,0.0,964.9,0,0,95635
4681,1,1,0,0,9,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,83.85,790.15,1,73,14,10.04,3723,1,Grizzly Flats,0,1,Cable,38.636102,-120.522149,0,87.204,0,0,None,659,0,1,0,0,9,2,111.0,90.36,0.0,790.15,0,0,95636
4682,0,1,0,0,27,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Credit card (automatic),88.3,2467.75,1,72,12,16.94,2420,1,Guinda,1,0,DSL,38.830739,-122.196202,0,91.83200000000001,0,0,None,228,0,0,0,0,27,0,296.0,457.38000000000005,0.0,2467.75,0,0,95637
4683,1,0,0,0,24,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.1,2322.85,0,60,14,30.42,3192,0,Herald,0,1,DSL,38.313447,-121.12388600000001,0,94.1,0,0,Offer C,1745,0,0,0,1,24,2,0.0,730.08,0.0,2322.85,0,1,95638
4684,1,0,0,0,69,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),104.05,7262,1,50,26,2.52,4254,1,Hood,1,1,Cable,38.375325,-121.507935,0,108.212,0,0,None,213,1,0,0,1,69,1,1888.0,173.88,0.0,7262.0,0,0,95639
4685,0,0,1,0,46,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),108.9,4854.3,0,29,48,2.0,5119,0,Ione,1,0,DSL,38.33788,-120.954202,1,108.9,0,6,None,9752,1,0,1,1,46,1,2330.0,92.0,0.0,4854.3,1,0,95640
4686,0,1,0,0,72,1,1,Fiber optic,1,1,0,1,Two year,1,Bank transfer (automatic),107.4,7748.75,0,66,18,31.31,5294,0,Isleton,1,0,Fiber Optic,38.154823,-121.601358,0,107.4,0,0,None,2010,1,0,0,1,72,0,0.0,2254.32,0.0,7748.75,0,1,95641
4687,1,0,1,0,22,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),94.7,1914.9,1,52,16,37.8,5615,1,Jackson,1,1,Fiber Optic,38.336216,-120.76901000000001,1,98.488,0,7,None,6202,0,0,1,1,22,3,0.0,831.5999999999998,0.0,1914.9,0,1,95642
4688,0,1,1,0,70,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,90.85,6470.1,0,68,25,38.5,5129,0,Knights Landing,0,0,DSL,38.875508,-121.76586599999999,1,90.85,0,10,None,1793,0,1,1,1,70,1,0.0,2695.0,0.0,6470.1,0,1,95645
4689,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.9,57.4,0,52,0,26.9,2822,0,Kirkwood,0,0,NA,38.631489,-120.01516699999999,0,19.9,0,0,Offer E,129,0,0,0,0,2,1,0.0,53.8,0.0,57.4,0,0,95646
4690,1,0,1,0,31,1,0,DSL,0,0,0,1,Month-to-month,1,Credit card (automatic),66.4,2019.8,0,56,28,25.3,3282,0,Lincoln,1,1,Fiber Optic,38.922812,-121.312005,1,66.4,0,7,Offer C,15286,1,0,1,1,31,1,0.0,784.3000000000002,0.0,2019.8,0,1,95648
4691,0,1,1,0,56,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),100.65,5688.05,1,68,32,33.81,4803,1,Loomis,1,0,Cable,38.809175,-121.171375,1,104.67600000000002,0,1,None,11191,0,0,1,0,56,4,0.0,1893.36,0.0,5688.05,0,1,95650
4692,0,0,1,1,16,1,0,Fiber optic,1,0,1,1,Month-to-month,0,Bank transfer (automatic),100.7,1522.7,0,57,76,27.27,3337,0,Lotus,1,0,Cable,38.815515000000005,-120.916997,1,100.7,3,10,Offer D,485,0,1,1,1,16,2,1157.0,436.32,0.0,1522.7,0,0,95651
4693,1,0,0,1,52,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.6,1334.5,0,26,0,23.12,5662,0,Madison,0,1,NA,38.674276,-121.96186599999999,0,25.6,1,0,None,844,0,0,0,0,52,2,0.0,1202.24,0.0,1334.5,1,0,95653
4694,1,0,1,1,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.85,252,0,35,0,40.2,2928,0,Mather,0,1,NA,38.549822,-121.266725,1,19.85,3,1,Offer D,929,0,0,1,0,13,2,0.0,522.6,0.0,252.0,0,0,95655
4695,0,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.75,700.45,0,34,0,35.5,4261,0,Newcastle,0,0,NA,38.883224,-121.15918,0,20.75,0,0,Offer C,6096,0,0,0,0,35,0,0.0,1242.5,0.0,700.45,0,0,95658
4696,0,0,0,0,59,1,0,Fiber optic,0,0,1,1,Two year,0,Electronic check,95.8,5655.45,0,36,30,30.44,5470,0,Nicolaus,1,0,Fiber Optic,38.788897999999996,-121.608624,0,95.8,0,0,None,751,0,0,0,1,59,0,1697.0,1795.96,0.0,5655.45,0,0,95659
4697,1,0,1,0,72,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.65,6747.35,0,39,23,33.22,5943,0,North Highlands,1,1,Fiber Optic,38.671295,-121.388251,1,94.65,0,9,None,32202,0,0,1,1,72,0,0.0,2391.84,0.0,6747.35,0,1,95660
4698,0,1,1,0,66,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),80.55,5265.1,1,74,3,21.7,4400,1,Roseville,1,0,Cable,38.736684999999994,-121.25198400000001,1,83.772,0,1,None,25173,0,0,1,0,66,2,158.0,1432.2,0.0,5265.1,0,0,95661
4699,0,0,1,0,49,1,1,Fiber optic,1,1,0,1,Two year,0,Credit card (automatic),106.65,5174.35,0,35,12,40.67,5948,0,Orangevale,1,0,Fiber Optic,38.689174,-121.21843500000001,1,106.65,0,10,None,32040,1,0,1,1,49,2,621.0,1992.83,0.0,5174.35,0,0,95662
4700,0,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.85,105.6,0,43,29,5.47,2245,0,Penryn,0,0,Fiber Optic,38.859093,-121.182872,0,45.85,0,0,Offer E,2048,0,2,0,0,2,1,31.0,10.94,0.0,105.6,0,0,95663
4701,1,1,0,0,21,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.35,2271.85,0,75,17,24.91,4934,0,Pilot Hill,1,1,Fiber Optic,38.803731,-121.04379899999999,0,104.35,0,0,Offer D,1173,0,0,0,1,21,1,386.0,523.11,0.0,2271.85,0,0,95664
4702,1,1,0,0,54,0,No phone service,DSL,0,1,1,1,One year,1,Electronic check,55.45,2966.95,0,72,26,0.0,4521,0,Pine Grove,1,1,Fiber Optic,38.400264,-120.641274,0,55.45,0,0,None,4354,0,0,0,1,54,1,0.0,0.0,0.0,2966.95,0,1,95665
4703,1,1,1,0,24,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,78.85,1772.25,1,71,24,2.05,3079,1,Pioneer,0,1,Fiber Optic,38.546999,-120.27111399999998,1,82.00399999999998,0,1,None,5501,0,1,1,0,24,4,425.0,49.2,0.0,1772.25,0,0,95666
4704,1,0,0,0,1,1,1,DSL,1,1,0,0,Month-to-month,0,Electronic check,61.15,61.15,0,47,3,17.07,4592,0,Placerville,0,1,Fiber Optic,38.733714,-120.79521299999999,0,61.15,0,0,Offer E,34146,0,0,0,0,1,2,0.0,17.07,0.0,61.15,0,0,95667
4705,1,0,0,0,6,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,78.95,494.95,0,55,28,29.52,4093,0,Pleasant Grove,0,1,DSL,38.833554,-121.498102,0,78.95,0,0,Offer E,901,0,0,0,0,6,0,0.0,177.12,0.0,494.95,0,1,95668
4706,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.45,44.45,1,63,24,48.31,4879,1,Plymouth,0,0,DSL,38.489273,-120.89161399999999,0,46.228,0,0,Offer E,2220,0,1,0,0,1,2,0.0,48.31,0.0,44.45,0,1,95669
4707,1,0,0,1,49,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),109.2,5290.45,0,35,58,4.76,6005,0,Rancho Cordova,1,1,Cable,38.602723,-121.279913,0,109.2,3,0,None,49729,0,0,0,1,49,0,3068.0,233.24,0.0,5290.45,0,0,95670
4708,0,0,1,1,56,1,0,DSL,1,1,0,0,Two year,1,Credit card (automatic),61.3,3346.8,0,59,53,18.99,4173,0,Rescue,1,0,Cable,38.724321999999994,-120.99123700000001,1,61.3,3,7,None,3815,0,0,1,0,56,1,0.0,1063.4399999999996,0.0,3346.8,0,1,95672
4709,0,1,0,0,56,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,96.85,5219.65,0,69,18,46.67,5679,0,Rio Linda,0,0,DSL,38.688764,-121.457596,0,96.85,0,0,None,14010,0,1,0,1,56,1,0.0,2613.52,0.0,5219.65,0,1,95673
4710,0,0,1,1,6,0,No phone service,DSL,0,1,0,0,Two year,0,Mailed check,40.55,217.5,0,61,10,0.0,2866,0,Rio Oso,1,0,DSL,38.954144,-121.48253600000001,1,40.55,2,7,Offer E,947,1,0,1,0,6,2,22.0,0.0,0.0,217.5,0,0,95674
4711,1,0,0,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.8,607.7,0,55,0,41.52,4636,0,River Pines,0,1,NA,38.545775,-120.743325,0,19.8,0,0,Offer C,364,0,0,0,0,32,1,0.0,1328.64,0.0,607.7,0,0,95675
4712,1,0,1,1,50,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,108.25,5431.4,0,34,19,41.58,4972,0,Rocklin,1,1,Fiber Optic,38.7904,-121.23697299999999,1,108.25,1,3,None,21510,0,0,1,1,50,0,1032.0,2079.0,0.0,5431.4,0,0,95677
4713,1,0,1,1,58,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),105.05,6004.85,0,33,10,33.82,5870,0,Roseville,1,1,Fiber Optic,38.759751,-121.288545,1,105.05,2,2,None,30614,1,0,1,1,58,1,0.0,1961.56,0.0,6004.85,0,1,95678
4714,0,0,1,1,65,1,1,DSL,1,1,1,1,Two year,1,Mailed check,90.45,5957.9,0,43,14,28.46,5509,0,Sheridan,1,0,Cable,38.984756,-121.345074,1,90.45,1,3,None,1219,1,0,1,1,65,0,834.0,1849.9,0.0,5957.9,0,0,95681
4715,0,0,0,0,64,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),86.4,5442.05,0,21,73,8.52,6474,0,Shingle Springs,1,0,Cable,38.598936,-120.96309199999999,0,86.4,0,0,None,24738,1,2,0,1,64,1,0.0,545.28,0.0,5442.05,1,1,95682
4716,0,0,1,0,66,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),66.9,4370.25,0,49,11,44.4,5546,0,Sloughhouse,1,0,Fiber Optic,38.470423,-121.114897,1,66.9,0,5,Offer A,4731,0,0,1,0,66,0,48.07,2930.4,0.0,4370.25,0,1,95683
4717,1,0,1,0,38,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,110.7,4428.6,0,59,15,42.08,5461,0,Somerset,1,1,Fiber Optic,38.606703,-120.58665900000001,1,110.7,0,9,Offer C,2958,1,0,1,1,38,2,66.43,1599.04,0.0,4428.6,0,1,95684
4718,0,0,1,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.0,416.45,0,21,0,19.15,3585,0,Sutter Creek,0,0,NA,38.432145,-120.77068999999999,1,20.0,0,2,Offer D,4610,0,0,1,0,20,1,0.0,383.0,0.0,416.45,1,0,95685
4719,1,0,0,0,36,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.9,3067.2,1,46,24,24.66,2455,1,Thornton,0,1,DSL,38.157794,-121.520223,0,88.296,0,0,None,1472,0,0,0,1,36,0,736.0,887.76,0.0,3067.2,0,0,95686
4720,1,1,0,0,64,1,1,Fiber optic,0,0,1,1,One year,0,Electronic check,102.1,6688.1,0,67,26,10.07,6100,0,Vacaville,1,1,Cable,38.333133000000004,-121.920151,0,102.1,0,0,None,63157,1,2,0,1,64,4,1739.0,644.48,0.0,6688.1,0,0,95687
4721,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.25,20.25,1,41,0,23.16,2959,1,Vacaville,0,1,NA,38.419088,-122.02456799999999,0,20.25,0,0,Offer E,32564,0,0,0,0,1,3,0.0,23.16,0.0,20.25,0,0,95688
4722,0,0,0,0,60,1,0,DSL,0,1,1,0,One year,1,Credit card (automatic),70.15,4224.7,0,49,2,38.88,4260,0,Volcano,1,0,DSL,38.481902000000005,-120.603668,0,70.15,0,0,None,1273,1,0,0,0,60,0,84.0,2332.8,0.0,4224.7,0,0,95689
4723,1,0,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.35,74.35,1,56,12,4.8,5633,1,Walnut Grove,0,1,Fiber Optic,38.240419,-121.587535,0,77.324,0,0,None,2344,0,0,0,0,1,2,0.0,4.8,0.0,74.35,0,0,95690
4724,0,0,1,1,50,1,1,DSL,1,1,0,1,One year,1,Bank transfer (automatic),80.05,4042.2,0,50,76,49.18,5823,0,West Sacramento,1,0,Cable,38.627951,-121.59328700000002,1,80.05,3,6,Offer B,19050,1,0,1,1,50,1,0.0,2459.0,0.0,4042.2,0,1,95691
4725,1,0,0,0,1,1,1,DSL,0,0,0,0,Month-to-month,0,Mailed check,62.05,62.05,1,58,13,47.83,2937,1,Wheatland,1,1,DSL,39.043387,-121.40983700000001,0,64.532,0,0,Offer E,3600,1,1,0,0,1,2,0.0,47.83,0.0,62.05,0,0,95692
4726,0,0,1,0,72,0,No phone service,DSL,1,1,0,1,Two year,1,Electronic check,49.2,3580.95,0,57,15,0.0,4700,0,Wilton,1,0,DSL,38.392559000000006,-121.22509299999999,1,49.2,0,2,Offer A,5889,0,0,1,1,72,1,537.0,0.0,0.0,3580.95,0,0,95693
4727,1,0,1,0,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.5,1198.8,0,28,0,31.29,5848,0,Winters,0,1,NA,38.578604,-122.024579,1,20.5,0,9,Offer B,8406,0,0,1,0,60,1,0.0,1877.4,0.0,1198.8,1,0,95694
4728,1,0,0,0,46,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,38.25,1755.35,0,40,2,0.0,2653,0,Woodland,1,1,Cable,38.71967,-121.862416,0,38.25,0,0,Offer B,38547,1,0,0,0,46,0,35.0,0.0,0.0,1755.35,0,0,95695
4729,0,0,1,1,69,0,No phone service,DSL,0,1,1,1,Two year,1,Credit card (automatic),54.95,3772.5,0,60,56,0.0,4175,0,Alta,1,0,Fiber Optic,39.218096,-120.79153000000001,1,54.95,3,4,Offer A,751,0,2,1,1,69,1,0.0,0.0,0.0,3772.5,0,1,95701
4730,1,1,0,0,31,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),96.6,2877.95,0,68,10,15.35,3364,0,Applegate,1,1,Cable,38.983388,-120.98881399999999,0,96.6,0,0,Offer C,1526,1,1,0,0,31,2,28.78,475.85,0.0,2877.95,0,1,95703
4731,1,0,1,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.9,357.7,0,49,0,32.47,5964,0,Camino,0,1,NA,38.748315999999996,-120.67551200000001,1,19.9,3,2,Offer D,4829,0,2,1,0,19,1,0.0,616.93,0.0,357.7,0,0,95709
4732,0,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.9,1397.3,0,28,0,20.49,6015,0,Colfax,0,0,NA,39.084645,-120.89401399999998,1,19.9,2,1,Offer A,8525,0,0,1,0,71,1,0.0,1454.79,0.0,1397.3,1,0,95713
4733,1,0,1,0,12,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,84.6,959.9,0,62,7,39.0,2499,0,Dutch Flat,1,1,DSL,39.197215,-120.83679,1,84.6,0,9,Offer D,350,0,0,1,0,12,1,0.0,468.0,0.0,959.9,0,1,95714
4734,1,0,1,1,39,1,0,DSL,1,0,1,1,One year,0,Credit card (automatic),80.0,3182.95,1,42,10,35.7,2704,1,Emigrant Gap,1,1,DSL,39.23754,-120.720196,1,83.2,0,1,None,185,1,0,1,1,39,0,318.0,1392.3000000000004,0.0,3182.95,0,0,95715
4735,1,0,0,0,44,1,1,DSL,0,1,1,1,One year,1,Bank transfer (automatic),85.25,3704.15,0,54,21,49.57,2292,0,Gold Run,1,1,Fiber Optic,39.170376,-120.838404,0,85.25,0,0,Offer B,407,1,0,0,1,44,0,0.0,2181.08,0.0,3704.15,0,1,95717
4736,0,0,1,1,56,1,1,DSL,1,1,1,0,Two year,0,Credit card (automatic),81.25,4620.4,0,51,30,25.9,5907,0,Kyburz,1,0,Fiber Optic,38.766036,-120.209673,1,81.25,2,10,Offer B,183,1,0,1,0,56,0,0.0,1450.4,0.0,4620.4,0,1,95720
4737,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),115.5,8312.75,0,26,76,24.32,4697,0,Echo Lake,1,0,Fiber Optic,38.851842,-120.076204,1,115.5,0,4,Offer A,69,1,0,1,1,72,0,6318.0,1751.04,0.0,8312.75,1,0,95721
4738,1,0,0,0,5,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Mailed check,104.1,541.9,1,43,9,38.89,3131,1,Meadow Vista,1,1,Fiber Optic,39.003358,-121.022539,0,108.264,0,0,Offer E,3747,0,0,0,1,5,0,49.0,194.45,0.0,541.9,0,0,95722
4739,0,0,0,0,11,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Bank transfer (automatic),79.0,929.3,0,28,48,10.06,3885,0,Pollock Pines,0,0,Cable,38.733908,-120.45341599999999,0,79.0,0,0,Offer D,8577,0,0,0,0,11,0,44.61,110.66,0.0,929.3,1,1,95726
4740,1,1,1,0,24,0,No phone service,DSL,1,0,0,1,Month-to-month,0,Bank transfer (automatic),39.1,971.3,1,75,6,0.0,4591,1,Soda Springs,0,1,Cable,39.279068,-120.414275,1,40.664,0,1,None,88,0,0,1,0,24,0,0.0,0.0,0.0,971.3,0,1,95728
4741,0,1,1,0,15,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,94.65,1285.05,0,66,19,37.84,5868,0,Twin Bridges,0,0,Cable,38.805481,-120.13287,1,94.65,0,5,Offer D,25,0,0,1,1,15,2,244.0,567.6,0.0,1285.05,0,0,95735
4742,1,0,0,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.8,1521.2,0,31,0,23.43,4626,0,Weimar,0,1,NA,39.00978,-120.978273,0,20.8,0,0,Offer A,31,0,0,0,0,72,1,0.0,1686.96,0.0,1521.2,0,0,95736
4743,1,0,1,0,56,1,1,DSL,0,1,0,0,Two year,0,Credit card (automatic),59.5,3389.25,0,34,17,35.55,5477,0,Rancho Cordova,1,1,Fiber Optic,38.591134000000004,-121.161585,1,59.5,0,9,Offer B,299,0,0,1,0,56,2,576.0,1990.8,0.0,3389.25,0,0,95742
4744,1,1,0,0,64,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.05,1198.05,0,79,0,4.99,4309,0,Granite Bay,0,1,NA,38.749466,-121.184196,0,20.05,0,0,None,20675,0,0,0,0,64,0,0.0,319.36,0.0,1198.05,0,0,95746
4745,0,0,1,0,34,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.45,3414.65,0,20,47,35.29,3744,0,Roseville,1,0,DSL,38.784329,-121.373245,1,100.45,0,10,Offer C,25418,0,0,1,1,34,1,0.0,1199.86,0.0,3414.65,1,1,95747
4746,1,0,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.5,162.45,1,30,33,17.22,5944,1,Elk Grove,0,1,Fiber Optic,38.353629999999995,-121.44195,0,79.56,0,0,Offer E,47065,0,0,0,0,2,4,0.0,34.44,0.0,162.45,0,1,95758
4747,1,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.6,754,0,22,0,42.02,2858,0,El Dorado Hills,0,1,NA,38.684437,-121.05563400000001,0,20.6,0,0,Offer C,22028,0,0,0,0,35,3,0.0,1470.7,0.0,754.0,1,0,95762
4748,1,0,0,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.3,467.15,0,24,0,23.03,2768,0,Rocklin,0,1,NA,38.823278,-121.281856,0,20.3,0,0,Offer D,15494,0,0,0,0,22,2,0.0,506.66,0.0,467.15,1,0,95765
4749,1,0,0,0,5,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.2,216.9,1,47,20,7.31,4336,1,Woodland,0,1,Fiber Optic,38.694081,-121.69443100000001,0,51.168000000000006,0,0,Offer E,15022,1,0,0,0,5,5,43.0,36.55,0.0,216.9,0,0,95776
4750,1,0,0,0,9,0,No phone service,DSL,1,1,0,0,One year,0,Mailed check,39.55,373,0,34,19,0.0,3755,0,Sacramento,1,1,Fiber Optic,38.584505,-121.491956,0,39.55,0,0,Offer E,16599,0,0,0,0,9,0,71.0,0.0,0.0,373.0,0,0,95814
4751,1,0,0,0,11,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),23.15,245.2,1,42,0,30.91,5671,1,Sacramento,0,1,NA,38.608405,-121.449942,0,23.15,0,0,None,25355,0,0,0,0,11,1,0.0,340.01,0.0,245.2,0,0,95815
4752,1,0,0,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.45,481.1,0,56,0,46.17,3434,0,Sacramento,0,1,NA,38.574856,-121.46503999999999,0,20.45,0,0,Offer D,16164,0,0,0,0,23,0,0.0,1061.91,0.0,481.1,0,0,95816
4753,0,0,1,1,4,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,80.85,302.75,1,22,65,44.28,2961,1,Sacramento,0,0,Cable,38.550722,-121.457314,1,84.084,0,1,Offer E,14966,0,1,1,1,4,2,197.0,177.12,0.0,302.75,1,0,95817
4754,1,0,1,0,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.25,1728.2,0,47,0,22.83,4571,0,Sacramento,0,1,NA,38.556306,-121.49581699999999,1,25.25,0,5,Offer A,21313,0,0,1,0,68,2,0.0,1552.4399999999996,0.0,1728.2,0,0,95818
4755,1,0,1,0,33,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,91.25,2964.05,0,55,17,26.8,3296,0,Sacramento,0,1,Fiber Optic,38.567594,-121.43750700000001,1,91.25,0,1,Offer C,15975,0,0,1,1,33,0,504.0,884.4,0.0,2964.05,0,0,95819
4756,1,0,0,0,31,1,0,DSL,1,1,1,0,Month-to-month,1,Bank transfer (automatic),72.45,2156.25,0,48,27,41.23,3175,0,Sacramento,1,1,DSL,38.53508,-121.444144,0,72.45,0,0,None,37031,1,0,0,0,31,2,582.0,1278.13,0.0,2156.25,0,0,95820
4757,1,0,0,0,1,1,1,DSL,0,1,0,0,Month-to-month,0,Mailed check,60.1,60.1,1,26,94,23.63,5654,1,Sacramento,0,1,DSL,38.625096,-121.38365800000001,0,62.50400000000001,0,0,Offer E,35426,1,3,0,0,1,3,0.0,23.63,0.0,60.1,1,0,95821
4758,0,0,0,0,56,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.7,1051.9,0,42,0,32.88,4831,0,Sacramento,0,0,NA,38.512569,-121.49518400000001,0,19.7,0,0,Offer B,44683,0,0,0,0,56,1,0.0,1841.28,0.0,1051.9,0,0,95822
4759,1,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,78.95,78.95,1,62,24,23.96,2038,1,Sacramento,0,1,Fiber Optic,38.475465,-121.443625,0,82.10799999999999,0,0,Offer E,72199,0,0,0,0,1,2,0.0,23.96,0.0,78.95,0,0,95823
4760,1,0,1,1,66,1,0,DSL,1,1,1,0,One year,1,Electronic check,75.1,5013,0,59,76,29.5,6123,0,Sacramento,1,1,Fiber Optic,38.517295000000004,-121.439819,1,75.1,3,0,Offer A,30580,1,0,0,0,66,2,380.99,1947.0,0.0,5013.0,0,1,95824
4761,1,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.0,1738.9,0,22,0,19.04,4275,0,Sacramento,0,1,NA,38.590035,-121.41245500000001,1,25.0,2,3,Offer A,30715,0,0,1,0,72,1,0.0,1370.88,0.0,1738.9,1,0,95825
4762,1,1,0,0,34,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),69.15,2275.1,0,67,30,13.56,4478,0,Sacramento,0,1,DSL,38.542532,-121.378826,0,69.15,0,0,Offer C,38818,0,0,0,0,34,2,683.0,461.04,0.0,2275.1,0,0,95826
4763,0,0,1,1,58,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,91.55,5511.65,0,49,17,40.74,6423,0,Sacramento,1,0,Fiber Optic,38.549184999999994,-121.32838600000001,1,91.55,2,5,Offer B,19611,0,0,1,0,58,1,0.0,2362.92,0.0,5511.65,0,1,95827
4764,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.15,98.5,1,56,23,6.47,2699,1,Sacramento,0,1,DSL,38.486938,-121.39580500000001,0,46.956,0,0,Offer E,54880,0,0,0,0,2,2,2.27,12.94,0.0,98.5,0,1,95828
4765,1,0,0,0,37,0,No phone service,DSL,0,0,1,0,Two year,0,Credit card (automatic),35.8,1316.9,0,51,25,0.0,5658,0,Sacramento,0,1,DSL,38.486502,-121.334051,0,35.8,0,0,None,11396,0,0,0,0,37,0,329.0,0.0,0.0,1316.9,0,0,95829
4766,0,0,0,0,71,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),113.15,7993.3,0,25,76,28.4,4955,0,Sacramento,1,0,Fiber Optic,38.490508,-121.284171,0,113.15,0,0,Offer A,592,1,0,0,1,71,0,0.0,2016.4,0.0,7993.3,1,1,95830
4767,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.85,19.85,0,55,0,47.46,2618,0,Sacramento,0,1,NA,38.494832,-121.52944699999999,1,19.85,1,5,None,42832,0,0,1,0,1,0,0.0,47.46,0.0,19.85,0,0,95831
4768,1,1,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.8,1388.45,0,77,0,32.12,5819,0,Sacramento,0,1,NA,38.445939,-121.49685500000001,1,19.8,1,5,None,9063,0,0,1,0,71,1,0.0,2280.52,0.0,1388.45,0,0,95832
4769,1,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.9,666,0,63,0,24.23,2334,0,Sacramento,0,1,NA,38.619049,-121.517552,1,19.9,2,7,None,31422,0,0,1,0,35,1,0.0,848.0500000000002,0.0,666.0,0,0,95833
4770,0,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.7,94.45,0,62,0,44.13,4122,0,Sacramento,0,0,NA,38.646209000000006,-121.52446,1,19.7,3,5,None,8403,0,0,1,0,6,1,0.0,264.78000000000003,0.0,94.45,0,0,95834
4771,0,0,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.4,244.65,1,28,84,46.6,2448,1,Sacramento,0,0,Cable,38.685069,-121.543709,0,82.57600000000002,0,0,Offer E,854,0,0,0,0,3,3,206.0,139.8,0.0,244.65,1,0,95835
4772,0,0,1,1,69,1,0,DSL,0,1,0,0,One year,0,Bank transfer (automatic),59.1,4134.7,0,47,19,14.48,5846,0,Sacramento,1,0,Cable,38.691607,-121.60228400000001,1,59.1,1,5,Offer A,264,1,0,1,0,69,0,786.0,999.12,0.0,4134.7,0,0,95837
4773,1,0,0,0,44,0,No phone service,DSL,0,1,1,1,One year,1,Mailed check,53.95,2375.4,1,38,4,0.0,3051,1,Sacramento,1,1,Fiber Optic,38.646096,-121.44243300000001,0,56.108,0,0,Offer B,34894,0,0,0,1,44,3,0.0,0.0,0.0,2375.4,0,1,95838
4774,0,0,1,0,53,1,1,Fiber optic,0,0,0,1,One year,1,Electronic check,91.15,4862.5,0,21,53,42.18,6439,0,Sacramento,0,0,Fiber Optic,38.660441999999996,-121.346321,1,91.15,0,2,Offer B,20993,1,0,1,1,53,1,0.0,2235.54,0.0,4862.5,1,1,95841
4775,0,0,1,0,24,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),99.3,2431.35,1,63,31,44.96,4811,1,Sacramento,1,0,Cable,38.687367,-121.34848000000001,1,103.272,0,0,None,31373,0,0,0,1,24,2,754.0,1079.04,0.0,2431.35,0,0,95842
4776,0,0,1,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,68.95,351.5,0,58,10,18.65,5536,0,Antelope,0,0,Fiber Optic,38.715498,-121.36341100000001,1,68.95,0,0,None,36432,0,0,0,0,5,2,0.0,93.25,0.0,351.5,0,1,95843
4777,0,0,0,1,2,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,51.55,106.2,0,21,27,18.61,4057,0,Sacramento,0,0,DSL,38.585826000000004,-121.376263,0,51.55,1,0,None,23362,0,0,0,0,2,1,29.0,37.22,0.0,106.2,1,0,95864
4778,1,0,0,1,62,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.4,1413,0,62,0,17.56,4889,0,Marysville,0,1,NA,39.19514,-121.503883,0,24.4,1,0,Offer B,38091,0,0,0,0,62,0,0.0,1088.72,0.0,1413.0,0,0,95901
4779,0,0,1,0,19,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.8,1743.05,0,58,23,10.68,3249,0,Beale Afb,1,0,Fiber Optic,39.125310999999996,-121.392283,1,96.8,0,9,Offer D,5654,0,0,1,1,19,0,0.0,202.92,0.0,1743.05,0,1,95903
4780,1,0,0,0,9,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.05,657.5,0,42,24,48.25,3522,0,Alleghany,0,1,DSL,39.467828000000004,-120.84138600000001,0,70.05,0,0,None,118,0,0,0,0,9,4,158.0,434.25,0.0,657.5,0,0,95910
4781,1,0,0,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.5,1050.5,0,29,0,24.17,5625,0,Arbuckle,0,1,NA,38.982372999999995,-122.047751,0,19.5,0,0,Offer B,4796,0,0,0,0,53,1,0.0,1281.01,0.0,1050.5,1,0,95912
4782,1,0,0,0,5,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Mailed check,78.75,426.35,0,32,24,32.91,2610,0,Bangor,0,1,Fiber Optic,39.396584999999995,-121.38028999999999,0,78.75,0,0,None,626,0,0,0,1,5,0,0.0,164.54999999999995,0.0,426.35,0,1,95914
4783,0,1,1,1,71,1,1,DSL,1,1,1,0,One year,0,Electronic check,69.2,4982.5,0,80,15,48.59,5546,0,Berry Creek,0,0,Fiber Optic,39.657228,-121.37778,1,69.2,1,7,None,1279,0,0,1,0,71,2,747.0,3449.890000000001,0.0,4982.5,0,0,95916
4784,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.55,19.55,0,44,0,10.2,5607,0,Biggs,0,0,NA,39.457388,-121.818201,0,19.55,0,0,None,3169,0,0,0,0,1,3,0.0,10.2,0.0,19.55,0,0,95917
4785,1,0,0,0,18,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.65,1451.9,1,58,8,38.87,3788,1,Browns Valley,0,1,Cable,39.292334000000004,-121.32059699999999,0,83.876,0,0,None,1477,0,0,0,0,18,0,116.0,699.66,0.0,1451.9,0,0,95918
4786,1,0,0,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,103.65,7634.8,0,64,16,10.87,6088,0,Brownsville,1,1,Fiber Optic,39.440687,-121.26358300000001,0,103.65,0,0,Offer A,1237,0,0,0,1,72,0,0.0,782.64,0.0,7634.8,0,1,95919
4787,0,0,1,0,4,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,54.7,235.05,0,36,3,6.77,3475,0,Butte City,0,0,Fiber Optic,39.449794,-121.93637199999999,1,54.7,0,2,None,303,0,0,1,0,4,1,7.0,27.08,0.0,235.05,0,0,95920
4788,1,0,0,0,59,1,1,DSL,0,0,0,0,Two year,0,Credit card (automatic),54.15,3116.15,0,35,9,49.48,4293,0,Camptonville,1,1,Fiber Optic,39.432127,-121.09928700000002,0,54.15,0,0,Offer B,632,0,1,0,0,59,1,28.05,2919.32,0.0,3116.15,0,1,95922
4789,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,71.1,71.1,1,41,10,10.19,5824,1,Canyon Dam,0,0,DSL,40.171312,-121.120605,0,73.944,0,0,Offer E,86,0,0,0,0,1,4,0.0,10.19,0.0,71.1,0,1,95923
4790,0,1,1,0,31,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.85,2633.4,0,68,3,5.3,5603,0,Challenge,0,0,DSL,39.461768,-121.195825,1,84.85,0,4,Offer C,262,0,0,1,1,31,0,79.0,164.29999999999995,0.0,2633.4,0,0,95925
4791,1,0,1,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.0,49.65,0,51,0,31.06,3985,0,Chico,0,1,NA,39.745712,-121.84333000000001,1,20.0,0,3,None,35808,0,0,1,0,3,0,0.0,93.18,0.0,49.65,0,0,95926
4792,0,1,1,0,65,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,106.25,6979.8,1,66,33,18.69,5965,1,Chico,1,0,DSL,39.681488,-121.83721000000001,1,110.5,0,1,None,32848,0,1,1,0,65,4,2303.0,1214.85,0.0,6979.8,0,0,95928
4793,1,0,1,0,49,1,0,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),99.25,4920.8,0,23,27,33.93,4995,0,Clipper Mills,1,1,Fiber Optic,39.562239,-121.14836000000001,1,99.25,0,4,Offer B,282,1,0,1,1,49,0,1329.0,1662.57,0.0,4920.8,1,0,95930
4794,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.35,46.35,0,42,0,44.34,5863,0,Colusa,0,1,NA,39.273096,-122.05076299999999,0,19.35,0,0,None,7503,0,0,0,0,2,0,0.0,88.68,0.0,46.35,0,0,95932
4795,0,0,1,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.8,1021.8,1,25,0,37.85,4166,1,Crescent Mills,0,0,NA,40.080342,-120.95780500000001,1,20.8,0,1,Offer B,178,0,0,1,0,53,0,0.0,2006.05,0.0,1021.8,1,0,95934
4796,0,0,1,0,55,1,0,Fiber optic,1,0,1,1,One year,1,Electronic check,94.75,5276.1,0,59,17,24.93,6021,0,Dobbins,0,0,DSL,39.381174,-121.21191,1,94.75,0,6,Offer B,614,0,0,1,1,55,2,0.0,1371.15,0.0,5276.1,0,1,95935
4797,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),114.05,8289.2,0,56,29,5.81,6254,0,Downieville,1,1,Fiber Optic,39.578792,-120.780786,1,114.05,1,4,Offer A,404,1,0,1,1,72,3,0.0,418.32,0.0,8289.2,0,1,95936
4798,0,1,0,0,36,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.9,2659.45,0,80,10,41.57,5041,0,Dunnigan,0,0,DSL,38.931425,-121.946081,0,74.9,0,0,Offer C,19,0,1,0,0,36,1,26.59,1496.52,0.0,2659.45,0,1,95937
4799,0,0,1,1,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),19.8,196.75,0,46,0,19.05,3196,0,Durham,0,0,NA,39.607831,-121.77795900000001,1,19.8,1,6,Offer D,3524,0,0,1,0,10,1,0.0,190.5,0.0,196.75,0,0,95938
4800,1,1,0,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.0,94,1,76,32,21.85,4176,1,Elk Creek,0,1,Cable,39.53222,-122.594879,0,97.76,0,0,None,587,0,0,0,0,1,0,0.0,21.85,0.0,94.0,0,0,95939
4801,0,0,1,1,72,1,1,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),80.85,5824.75,0,40,15,9.72,6317,0,Forbestown,1,0,Cable,39.531028000000006,-121.24807,1,80.85,2,5,Offer A,452,1,0,1,1,72,4,0.0,699.84,0.0,5824.75,0,1,95941
4802,0,0,0,0,28,1,0,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),54.65,1517.5,0,55,7,25.59,3185,0,Forest Ranch,0,0,DSL,40.077028000000006,-121.49416799999999,0,54.65,0,0,None,1351,1,0,0,0,28,0,106.0,716.52,0.0,1517.5,0,0,95942
4803,1,0,1,0,38,1,1,Fiber optic,1,0,1,0,Month-to-month,0,Bank transfer (automatic),91.7,3479.05,0,36,9,12.71,3676,0,Glenn,0,1,Fiber Optic,39.597975,-122.032248,1,91.7,0,3,None,1454,0,0,1,0,38,0,313.0,482.98,0.0,3479.05,0,0,95943
4804,0,0,0,0,61,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,118.6,7365.7,0,25,42,38.78,5536,0,Goodyears Bar,1,0,DSL,39.564113,-120.86883600000002,0,118.6,0,0,Offer B,76,1,0,0,1,61,2,3094.0,2365.58,0.0,7365.7,1,0,95944
4805,1,0,1,1,52,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.55,1331.05,0,34,0,29.55,5535,0,Grass Valley,0,1,NA,39.194539,-120.98806599999999,1,24.55,1,6,Offer B,23990,0,0,1,0,52,1,0.0,1536.6,0.0,1331.05,0,0,95945
4806,1,0,0,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.45,1195.95,0,45,0,9.05,5343,0,Penn Valley,0,1,NA,39.203817,-121.19583999999999,0,19.45,0,0,Offer A,9752,0,0,0,0,67,0,0.0,606.35,0.0,1195.95,0,0,95946
4807,0,0,0,1,34,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),116.15,3946.9,0,26,51,27.47,5104,0,Greenville,1,0,DSL,40.160385999999995,-120.83542800000001,0,116.15,3,0,None,2064,1,0,0,1,34,1,0.0,933.98,0.0,3946.9,1,1,95947
4808,0,0,0,0,54,1,0,DSL,1,0,1,1,Two year,0,Electronic check,80.6,4299.95,0,46,28,36.68,4231,0,Gridley,1,0,Fiber Optic,39.346897999999996,-121.75953700000001,0,80.6,0,0,None,9763,1,0,0,1,54,0,1204.0,1980.72,0.0,4299.95,0,0,95948
4809,0,0,1,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.3,20.3,0,60,0,6.64,4215,0,Grass Valley,0,0,NA,39.099204,-121.13796200000002,1,20.3,0,7,None,17922,0,0,1,0,1,0,0.0,6.64,0.0,20.3,0,0,95949
4810,0,1,0,0,15,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,89.85,1424.95,1,67,7,4.28,2668,1,Grimes,0,0,Cable,39.033058000000004,-121.89571799999999,0,93.444,0,0,Offer D,531,0,1,0,0,15,3,100.0,64.2,0.0,1424.95,0,0,95950
4811,0,0,0,0,4,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,46.0,193.6,1,48,18,15.07,5246,1,Hamilton City,0,0,DSL,39.732766999999996,-122.042298,0,47.84,0,0,None,1931,0,0,0,0,4,3,0.0,60.28,0.0,193.6,0,1,95951
4812,0,0,0,0,9,1,0,DSL,0,1,1,0,Month-to-month,0,Mailed check,66.25,620.55,1,27,76,24.81,5515,1,Live Oak,0,0,Cable,39.258746,-121.77696999999999,0,68.9,0,0,None,8695,1,3,0,0,9,3,472.0,223.29,0.0,620.55,1,0,95953
4813,0,0,0,1,46,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.8,4391.25,0,26,85,17.51,2405,0,Magalia,1,0,DSL,39.933852,-121.58437099999999,0,99.8,2,0,None,11168,0,0,0,1,46,1,0.0,805.46,0.0,4391.25,1,1,95954
4814,0,0,0,0,22,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,90.0,1993.8,1,60,25,12.19,4739,1,Maxwell,0,0,Cable,39.281194,-122.226568,0,93.6,0,0,None,1146,1,0,0,0,22,3,0.0,268.18,0.0,1993.8,0,1,95955
4815,1,0,0,0,38,1,0,Fiber optic,0,0,0,0,One year,1,Bank transfer (automatic),70.45,2597.6,1,39,19,33.71,5437,1,Meadow Valley,0,1,Cable,39.937017,-121.058043,0,73.268,0,0,None,301,0,1,0,0,38,1,494.0,1280.98,0.0,2597.6,0,0,95956
4816,0,0,1,1,55,1,1,DSL,1,1,1,0,One year,1,Credit card (automatic),75.0,4213.9,0,27,51,33.5,5011,0,Meridian,0,0,DSL,39.068071,-121.83263799999999,1,75.0,2,7,None,776,1,0,1,0,55,2,2149.0,1842.5,0.0,4213.9,1,0,95957
4817,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,19.9,0,21,0,1.5,5057,0,Nevada City,0,0,NA,39.333737,-120.858667,0,19.9,0,0,None,17269,0,0,0,0,1,1,0.0,1.5,0.0,19.9,1,0,95959
4818,1,1,1,0,64,1,0,Fiber optic,1,0,0,0,One year,0,Credit card (automatic),80.3,5017.7,0,77,16,14.87,4270,0,North San Juan,1,1,DSL,39.423046,-120.984472,1,80.3,0,5,None,565,0,0,1,0,64,0,803.0,951.68,0.0,5017.7,0,0,95960
4819,1,0,0,1,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.75,1052.35,1,62,0,26.21,6265,1,Olivehurst,0,1,NA,39.082568,-121.55325,0,19.75,0,0,Offer B,6439,0,0,0,0,53,3,0.0,1389.13,0.0,1052.35,0,0,95961
4820,0,0,1,0,58,1,1,DSL,1,0,1,1,Two year,1,Electronic check,84.3,4916.4,0,29,59,31.27,5724,0,Oregon House,1,0,Fiber Optic,39.342587,-121.24983300000001,1,84.3,0,1,None,1519,1,0,1,1,58,1,290.07,1813.66,0.0,4916.4,1,1,95962
4821,1,0,1,0,56,0,No phone service,DSL,0,0,1,1,One year,1,Bank transfer (automatic),54.05,2959.8,0,20,30,0.0,6445,0,Orland,1,1,Fiber Optic,39.748037,-122.30216899999999,1,54.05,0,10,None,13706,1,0,1,1,56,0,88.79,0.0,0.0,2959.8,1,1,95963
4822,1,0,1,1,72,1,0,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),104.9,7559.55,0,43,57,6.95,5169,0,Oroville,1,1,Fiber Optic,39.624561,-121.552866,1,104.9,3,5,Offer A,17782,1,0,1,1,72,2,4309.0,500.4,0.0,7559.55,0,0,95965
4823,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,53.95,53.95,1,49,12,31.16,2771,1,Oroville,0,1,Cable,39.473896,-121.415927,0,56.108,0,0,None,28382,1,0,0,0,1,5,0.0,31.16,0.0,53.95,0,1,95966
4824,1,1,1,0,72,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),97.25,7133.1,0,75,20,11.23,6156,0,Palermo,0,1,Cable,39.435756,-121.552071,1,97.25,0,7,None,1254,0,0,1,1,72,3,1427.0,808.5600000000002,0.0,7133.1,0,0,95968
4825,1,0,0,0,22,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,83.05,1799.3,0,35,16,11.46,5357,0,Paradise,0,1,Cable,39.69676,-121.644379,0,83.05,0,0,Offer D,28318,0,0,0,1,22,1,288.0,252.12,0.0,1799.3,0,0,95969
4826,0,1,0,0,8,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.5,829.55,1,79,16,45.16,5546,1,Princeton,1,0,Cable,39.424957,-122.03930700000001,0,109.72,0,0,None,495,0,0,0,0,8,4,133.0,361.28,0.0,829.55,0,0,95970
4827,0,0,0,1,16,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,81.0,1312.15,1,40,13,12.92,2335,1,Quincy,0,0,DSL,39.971228,-121.04116599999999,0,84.24000000000002,0,0,None,6189,0,1,0,0,16,1,171.0,206.72,0.0,1312.15,0,0,95971
4828,0,0,0,0,39,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Bank transfer (automatic),41.1,1597.05,0,35,8,0.0,3618,0,Chico,1,0,Fiber Optic,39.903271999999994,-121.843567,0,41.1,0,0,None,26971,1,0,0,0,39,2,12.78,0.0,0.0,1597.05,0,1,95973
4829,0,0,0,0,12,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),45.0,524.35,0,47,13,36.11,4998,0,Richvale,0,0,Fiber Optic,39.495768,-121.747472,0,45.0,0,0,None,74,0,0,0,0,12,1,68.0,433.32,0.0,524.35,0,0,95974
4830,1,0,1,0,54,1,0,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),74.55,4191.45,0,48,25,14.18,4544,0,Rough And Ready,0,1,Fiber Optic,39.225634,-121.15616299999999,1,74.55,0,8,None,1601,0,0,1,1,54,0,1048.0,765.72,0.0,4191.45,0,0,95975
4831,0,0,0,0,18,0,No phone service,DSL,1,1,0,0,One year,1,Mailed check,40.2,711.95,0,28,48,0.0,4624,0,Smartville,0,0,DSL,39.176595,-121.291692,0,40.2,0,0,None,963,1,2,0,0,18,2,0.0,0.0,0.0,711.95,1,1,95977
4832,1,0,1,0,32,1,0,DSL,1,1,0,1,One year,0,Mailed check,70.5,2201.75,0,47,6,44.45,5870,0,Stirling City,0,1,Fiber Optic,39.904002,-121.527823,1,70.5,0,7,None,28,1,0,1,1,32,0,0.0,1422.4,0.0,2201.75,0,1,95978
4833,0,0,0,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.75,806.95,0,40,0,37.46,5678,0,Stonyford,0,0,NA,39.288127,-122.41584099999999,0,19.75,0,0,None,844,0,1,0,0,41,1,0.0,1535.86,0.0,806.95,0,0,95979
4834,1,0,1,1,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.65,1620.45,0,60,0,14.41,4444,0,Strawberry Valley,0,1,NA,39.584579999999995,-121.09325600000001,1,24.65,2,6,None,101,0,0,1,0,67,1,0.0,965.47,0.0,1620.45,0,0,95981
4835,1,0,1,0,65,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,104.25,6812.95,0,48,10,41.2,5089,0,Sutter,1,1,Fiber Optic,39.172777,-121.80584499999999,1,104.25,0,4,None,3193,0,0,1,1,65,1,0.0,2678.0,0.0,6812.95,0,1,95982
4836,0,0,0,0,25,1,1,DSL,1,1,1,0,Month-to-month,1,Bank transfer (automatic),78.35,1837.9,0,19,85,28.05,4855,0,Taylorsville,1,0,Fiber Optic,40.053684000000004,-120.74311599999999,0,78.35,0,0,None,513,1,0,0,0,25,1,0.0,701.25,0.0,1837.9,1,1,95983
4837,0,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.8,69.8,1,34,14,11.08,2123,1,Twain,0,0,Cable,40.022184,-121.06238400000001,1,72.592,0,1,None,73,0,1,1,0,1,3,0.0,11.08,0.0,69.8,0,1,95984
4838,0,0,1,0,67,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),109.7,7344.45,0,50,23,17.72,4017,0,Washington,1,0,Fiber Optic,39.34128,-120.78686699999999,1,109.7,0,6,None,145,1,0,1,1,67,1,0.0,1187.24,0.0,7344.45,0,1,95986
4839,1,1,0,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,73.75,545.15,1,78,8,32.4,5638,1,Williams,0,1,Cable,39.117537,-122.284654,0,76.7,0,0,None,4579,0,0,0,0,7,4,4.36,226.8,0.0,545.15,0,1,95987
4840,0,1,0,0,43,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Credit card (automatic),33.45,1500.25,0,73,18,0.0,4757,0,Willows,0,0,Fiber Optic,39.493990999999994,-122.286363,0,33.45,0,0,None,8812,0,0,0,0,43,0,0.0,0.0,0.0,1500.25,0,1,95988
4841,0,0,0,0,24,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,94.6,2283.15,0,37,3,35.56,3667,0,Yuba City,0,0,DSL,39.027409999999996,-121.61498200000001,0,94.6,0,0,None,34967,0,0,0,1,24,0,0.0,853.44,0.0,2283.15,0,1,95991
4842,1,1,0,0,9,1,1,DSL,1,0,0,0,Month-to-month,0,Electronic check,54.55,494.05,1,79,8,2.45,4656,1,Yuba City,0,1,Cable,39.075694,-121.70606000000001,0,56.732,0,0,Offer E,27786,0,0,0,0,9,0,40.0,22.05,0.0,494.05,0,0,95993
4843,1,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.2,1376.5,0,29,0,23.55,5463,0,Redding,0,1,NA,40.587919,-122.46473200000001,1,20.2,1,2,None,31586,0,0,1,0,69,3,0.0,1624.95,0.0,1376.5,1,0,96001
4844,0,0,0,1,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.3,755.4,0,28,0,10.23,4186,0,Redding,0,0,NA,40.527834000000006,-122.318749,0,20.3,3,0,None,30338,0,0,0,0,37,0,0.0,378.51,0.0,755.4,1,0,96002
4845,1,0,1,1,20,0,No phone service,DSL,1,0,0,0,Two year,1,Credit card (automatic),39.4,825.4,0,33,22,0.0,3899,0,Redding,1,1,Fiber Optic,40.677649,-122.29467,1,39.4,1,4,None,41476,1,0,1,0,20,0,0.0,0.0,0.0,825.4,0,1,96003
4846,1,0,0,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),69.15,488.65,0,54,7,21.12,4320,0,Adin,0,1,Fiber Optic,41.171578000000004,-120.91316100000002,0,69.15,0,0,None,615,0,0,0,0,7,2,34.0,147.84,0.0,488.65,0,0,96006
4847,0,1,0,0,37,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.25,2841.55,1,78,19,26.95,5859,1,Anderson,0,0,Fiber Optic,40.448632,-122.306657,0,79.3,0,0,Offer C,21418,0,1,0,0,37,4,53.99,997.15,0.0,2841.55,0,1,96007
4848,0,0,0,0,5,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,93.9,486.85,1,44,11,46.45,5435,1,Bella Vista,0,0,Cable,40.722733000000005,-122.10966599999999,0,97.656,0,0,None,899,0,0,0,1,5,1,0.0,232.25,0.0,486.85,0,1,96008
4849,1,0,0,0,41,0,No phone service,DSL,0,0,1,1,One year,1,Electronic check,51.35,2075.1,0,50,8,0.0,5622,0,Bieber,1,1,Cable,41.083464,-121.107929,0,51.35,0,0,None,595,0,0,0,1,41,0,0.0,0.0,0.0,2075.1,0,1,96009
4850,0,0,0,0,54,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),100.05,5299.65,0,36,20,34.27,4478,0,Big Bar,0,0,DSL,40.775271999999994,-123.28741399999998,0,100.05,0,0,None,269,0,0,0,1,54,2,1060.0,1850.58,0.0,5299.65,0,0,96010
4851,0,1,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.4,204.7,1,71,3,2.26,2491,1,Big Bend,0,0,Cable,41.096569,-121.87908200000001,0,73.21600000000002,0,0,Offer E,265,0,0,0,0,3,6,6.0,6.7799999999999985,0.0,204.7,0,0,96011
4852,1,1,0,0,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.3,1356.3,0,67,0,20.62,4042,0,Burney,0,1,NA,40.946785,-121.719489,0,20.3,0,0,None,4552,0,0,0,0,69,0,0.0,1422.78,0.0,1356.3,0,0,96013
4853,0,0,0,0,53,1,0,Fiber optic,0,1,0,1,One year,1,Credit card (automatic),94.45,5042.75,0,59,6,33.88,5452,0,Callahan,1,0,Cable,41.388397,-122.79463600000001,0,94.45,0,0,None,290,1,0,0,1,53,0,303.0,1795.64,0.0,5042.75,0,0,96014
4854,1,0,1,1,18,0,No phone service,DSL,0,1,1,0,One year,0,Credit card (automatic),46.4,812.4,0,25,59,0.0,4003,0,Canby,1,1,Fiber Optic,41.486953,-120.913975,1,46.4,2,2,None,417,0,0,1,0,18,1,47.93,0.0,0.0,812.4,1,1,96015
4855,1,0,1,0,64,1,0,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),104.05,6605.55,0,61,8,4.76,4337,0,Cassel,0,1,DSL,40.936285,-121.57269199999999,1,104.05,0,1,None,344,1,0,1,1,64,0,528.0,304.64,0.0,6605.55,0,0,96016
4856,0,0,1,1,31,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,91.15,2995.45,1,39,14,38.67,5219,1,Castella,0,0,Cable,41.121108,-122.33661299999999,1,94.796,0,1,None,228,0,2,1,1,31,4,419.0,1198.77,0.0,2995.45,0,0,96017
4857,0,0,0,0,20,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),24.9,505.95,0,41,21,0.0,5942,0,Shasta Lake,0,0,DSL,40.692523,-122.369876,0,24.9,0,0,None,6277,0,0,0,0,20,0,0.0,0.0,0.0,505.95,0,1,96019
4858,1,0,1,1,57,1,0,DSL,1,1,0,0,One year,0,Mailed check,59.6,3509.4,0,37,58,14.55,4778,0,Chester,0,1,DSL,40.243494,-121.15473300000001,1,59.6,3,7,None,2664,1,1,1,0,57,1,2035.0,829.35,0.0,3509.4,0,0,96020
4859,1,1,1,0,63,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),108.5,6991.9,0,73,18,37.12,6453,0,Corning,1,1,Fiber Optic,39.913777,-122.289984,1,108.5,0,1,None,13840,0,0,1,1,63,0,0.0,2338.56,0.0,6991.9,0,1,96021
4860,1,0,1,1,13,0,No phone service,DSL,1,1,0,0,Two year,0,Mailed check,40.55,590.35,0,58,57,0.0,2898,0,Cottonwood,0,1,Fiber Optic,40.336392,-122.44853300000001,1,40.55,3,0,None,12348,1,0,0,0,13,1,336.0,0.0,0.0,590.35,0,0,96022
4861,0,1,1,0,48,1,0,DSL,0,1,0,1,One year,1,Bank transfer (automatic),58.95,2789.7,0,65,2,34.43,4815,0,Dorris,0,0,Fiber Optic,41.949216,-122.05006200000001,1,58.95,0,10,None,1162,0,1,1,1,48,1,0.0,1652.64,0.0,2789.7,0,1,96023
4862,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.95,137.95,1,45,29,15.33,5390,1,Douglas City,0,0,Cable,40.586588,-122.903677,0,73.78800000000003,0,0,None,960,0,2,0,0,2,3,40.0,30.66,0.0,137.95,0,0,96024
4863,1,0,1,1,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.75,1123.15,0,60,0,29.64,4937,0,Dunsmuir,0,1,NA,41.212695000000004,-122.392067,1,20.75,2,8,None,2602,0,0,1,0,57,1,0.0,1689.48,0.0,1123.15,0,0,96025
4864,1,0,1,0,71,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),113.15,7953.25,0,50,3,27.16,4068,0,Etna,1,1,DSL,41.405193,-123.008567,1,113.15,0,8,None,2156,1,0,1,1,71,0,239.0,1928.36,0.0,7953.25,0,0,96027
4865,0,0,1,1,7,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,48.8,349.8,0,56,28,9.1,4785,0,Fall River Mills,0,0,Cable,41.017282,-121.46894499999999,1,48.8,2,1,Offer E,1902,0,0,1,0,7,0,98.0,63.7,0.0,349.8,0,0,96028
4866,0,0,0,0,16,1,1,DSL,0,0,0,1,Month-to-month,1,Bank transfer (automatic),63.05,1067.05,0,56,23,42.73,3214,0,Flournoy,0,0,Cable,39.847840000000005,-122.544556,0,63.05,0,0,None,84,0,0,0,1,16,1,245.0,683.68,0.0,1067.05,0,0,96029
4867,1,0,1,0,34,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,100.85,3527.3,0,21,41,33.55,5891,0,Forks Of Salmon,1,1,Fiber Optic,41.232128,-123.194748,1,100.85,0,8,None,170,0,0,1,1,34,0,0.0,1140.6999999999996,0.0,3527.3,1,1,96031
4868,0,0,1,0,37,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.5,3762,1,26,30,36.29,4233,1,Escondido,1,0,Cable,33.141265000000004,-116.967221,1,103.48,0,1,None,48690,0,1,1,1,37,2,1129.0,1342.73,0.0,3762.0,1,0,92027
4869,1,0,0,0,16,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,80.55,1248.9,0,58,8,34.18,5183,0,French Gulch,0,1,Fiber Optic,40.740138,-122.587476,0,80.55,0,0,None,373,0,0,0,0,16,0,100.0,546.88,0.0,1248.9,0,0,96033
4870,1,0,0,1,48,1,1,DSL,1,1,0,0,One year,1,Bank transfer (automatic),64.4,3035.35,0,39,53,26.24,2545,0,Gazelle,1,1,DSL,41.411315,-122.697236,0,64.4,3,0,None,392,0,0,0,0,48,0,0.0,1259.52,0.0,3035.35,0,1,96034
4871,1,0,1,1,58,1,0,DSL,0,1,1,1,One year,1,Credit card (automatic),75.2,4300.8,0,54,29,35.35,4559,0,Gerber,0,1,Cable,40.031940000000006,-122.176023,1,75.2,2,9,None,3357,1,0,1,1,58,1,0.0,2050.3,0.0,4300.8,0,1,96035
4872,0,0,1,0,72,1,1,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),84.9,6065.3,0,36,19,1.34,4447,0,Greenview,1,0,Fiber Optic,41.528541,-122.955018,1,84.9,0,7,None,295,1,0,1,1,72,0,1152.0,96.48,0.0,6065.3,0,0,96037
4873,0,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.3,144.95,0,51,0,7.32,4764,0,Grenada,0,0,NA,41.599978,-122.539381,0,19.3,0,0,None,616,0,0,0,0,7,2,0.0,51.24,0.0,144.95,0,0,96038
4874,0,0,0,0,38,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),83.9,3233.6,1,26,53,36.18,2157,1,Happy Camp,1,0,Fiber Optic,41.831901,-123.487478,0,87.25600000000001,0,0,None,1294,0,0,0,1,38,1,0.0,1374.84,0.0,3233.6,1,1,96039
4875,0,1,1,0,48,1,1,Fiber optic,1,1,1,1,Month-to-month,0,Electronic check,117.45,5438.9,1,76,6,43.04,5915,1,Hat Creek,1,0,Fiber Optic,40.789799,-121.474529,1,122.148,0,9,None,397,1,3,1,0,48,6,326.0,2065.92,0.0,5438.9,0,0,96040
4876,1,0,0,0,10,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,104.4,1081.45,1,37,2,8.38,5035,1,Fallbrook,1,1,Cable,33.362575,-117.299644,0,108.576,0,0,None,42239,0,0,0,1,10,0,2.16,83.80000000000003,0.0,1081.45,0,1,92028
4877,0,0,0,0,30,1,0,DSL,1,1,1,0,One year,0,Credit card (automatic),74.65,2308.6,0,52,13,4.22,5616,0,Hornbrook,1,0,Fiber Optic,41.962127,-122.52769599999999,0,74.65,0,0,None,1026,1,0,0,0,30,0,300.0,126.6,0.0,2308.6,0,0,96044
4878,1,0,1,0,31,1,1,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),59.05,1882.8,0,33,21,28.72,5841,0,Hyampom,0,1,DSL,40.648024,-123.465088,1,59.05,0,0,None,268,0,0,0,0,31,1,39.54,890.3199999999998,0.0,1882.8,0,1,96046
4879,0,1,0,0,46,1,1,DSL,0,0,0,1,One year,1,Credit card (automatic),69.1,3255.35,0,65,26,16.04,3856,0,Igo,1,0,DSL,40.524535,-122.647172,0,69.1,0,0,None,911,1,0,0,1,46,1,846.0,737.8399999999998,0.0,3255.35,0,0,96047
4880,1,0,1,0,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.55,1067.65,0,32,0,46.91,4745,0,Junction City,0,1,NA,40.913191999999995,-123.06597,1,20.55,0,4,None,734,0,1,1,0,50,1,0.0,2345.5,0.0,1067.65,0,0,96048
4881,1,0,1,0,28,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),76.55,2065.4,0,31,5,21.91,2085,0,Klamath River,0,1,DSL,41.816595,-122.94828700000001,1,76.55,0,10,None,482,1,0,1,0,28,1,0.0,613.48,0.0,2065.4,0,1,96050
4882,0,0,0,0,66,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),62.5,4136.4,0,52,15,0.0,4165,0,Lakehead,1,0,Fiber Optic,40.883853,-122.41825800000001,0,62.5,0,0,None,1236,1,0,0,1,66,1,620.0,0.0,0.0,4136.4,0,0,96051
4883,1,1,0,0,8,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,29.4,221.9,1,65,4,0.0,5971,1,Lewiston,1,1,DSL,40.704293,-122.803899,0,30.576,0,0,Offer E,1845,0,2,0,0,8,1,9.0,0.0,0.0,221.9,0,0,96052
4884,0,0,1,1,41,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),94.9,3848,0,25,59,43.19,3539,0,Lookout,1,0,DSL,41.280478,-121.160249,1,94.9,3,2,None,386,0,0,1,1,41,2,2270.0,1770.79,0.0,3848.0,1,0,96054
4885,1,1,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),111.65,8022.85,0,72,19,16.92,4406,0,Los Molinos,1,1,Fiber Optic,40.059385,-122.091481,1,111.65,0,4,None,3756,1,0,1,1,72,0,1524.0,1218.2400000000002,0.0,8022.85,0,0,96055
4886,0,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.9,173.15,0,29,0,16.2,2750,0,Mcarthur,0,0,NA,41.108309999999996,-121.36036200000001,0,19.9,0,0,Offer E,1554,0,1,0,0,7,1,0.0,113.4,0.0,173.15,1,0,96056
4887,0,0,1,1,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.45,781.25,0,26,0,2.86,5587,0,Mccloud,0,0,NA,41.251321999999995,-122.105209,1,20.45,2,6,None,1586,0,0,1,0,38,0,0.0,108.68,0.0,781.25,1,0,96057
4888,1,0,0,0,44,1,0,Fiber optic,1,1,1,1,One year,1,Electronic check,106.05,4510.8,0,25,41,38.33,4588,0,Macdoel,1,1,DSL,41.769709000000006,-121.92063,0,106.05,0,0,None,816,0,0,0,1,44,0,0.0,1686.52,0.0,4510.8,1,1,96058
4889,1,0,1,1,47,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),113.45,5317.8,0,58,19,9.19,3729,0,Manton,1,1,Fiber Optic,40.426679,-121.850421,1,113.45,1,7,None,598,1,0,1,1,47,0,0.0,431.93,0.0,5317.8,0,1,96059
4890,1,0,1,1,53,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,92.55,4779.45,0,25,52,24.33,4700,0,Mill Creek,0,1,Fiber Optic,40.331975,-121.460674,1,92.55,2,5,None,78,1,0,1,0,53,0,0.0,1289.49,0.0,4779.45,1,1,96061
4891,1,0,1,0,4,1,1,DSL,0,0,1,0,Month-to-month,0,Electronic check,65.6,250.1,0,49,3,10.13,4552,0,Millville,1,1,DSL,40.531257000000004,-122.14813899999999,1,65.6,0,7,Offer E,830,0,0,1,0,4,0,8.0,40.52,0.0,250.1,0,0,96062
4892,1,1,0,0,20,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.35,1745.2,0,78,9,25.51,4915,0,Mineral,0,1,DSL,40.408796,-121.579609,0,84.35,0,0,Offer D,124,0,0,0,0,20,1,0.0,510.2000000000001,0.0,1745.2,0,1,96063
4893,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.65,74.9,1,46,12,24.9,4655,1,Fallbrook,0,1,Fiber Optic,33.362575,-117.299644,0,46.43600000000001,0,0,None,42239,0,0,0,0,2,2,9.0,49.8,0.0,74.9,0,0,92028
4894,1,1,1,0,57,1,1,DSL,0,1,1,0,One year,1,Credit card (automatic),71.1,4140.1,0,72,10,48.16,5462,0,Montgomery Creek,1,1,Cable,40.877552,-121.885884,1,71.1,0,2,None,431,0,0,1,0,57,0,0.0,2745.12,0.0,4140.1,0,1,96065
4895,0,1,1,0,44,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,85.15,3670.5,0,70,6,44.44,2672,0,Mount Shasta,0,0,Fiber Optic,41.33832,-122.290756,1,85.15,0,4,None,7309,1,0,1,0,44,2,22.02,1955.36,0.0,3670.5,0,1,96067
4896,1,0,0,0,24,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,49.7,1167.8,0,25,73,38.68,5832,0,Nubieber,1,1,Fiber Optic,41.082471999999996,-121.19521499999999,0,49.7,0,0,None,240,0,0,0,0,24,0,852.0,928.32,0.0,1167.8,1,0,96068
4897,1,0,1,1,15,0,No phone service,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),30.2,469.65,0,59,16,0.0,5825,0,Oak Run,0,1,Fiber Optic,40.689243,-122.037023,1,30.2,2,8,None,829,0,0,1,0,15,1,75.0,0.0,0.0,469.65,0,0,96069
4898,0,0,0,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,25.25,58.9,1,62,30,0.0,2088,1,Old Station,0,0,DSL,40.656287,-121.42896499999999,0,26.26,0,0,None,182,0,1,0,0,3,3,18.0,0.0,0.0,58.9,0,0,96071
4899,0,0,0,1,4,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),84.05,333.55,1,21,76,41.72,5552,1,Palo Cedro,1,0,Cable,40.582399,-122.19551200000001,0,87.412,0,0,None,4931,0,1,0,1,4,2,253.0,166.88,0.0,333.55,1,0,96073
4900,1,1,1,0,37,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.7,3171.15,1,75,29,46.61,4712,1,Paskenta,0,1,Fiber Optic,39.884395,-122.58751299999999,1,89.12799999999999,0,1,Offer C,263,0,0,1,0,37,0,0.0,1724.57,0.0,3171.15,0,1,96074
4901,0,0,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.7,74.7,1,23,76,44.11,4692,1,Paynes Creek,0,0,Cable,40.343213,-121.81541200000001,0,77.688,0,0,Offer E,433,0,1,0,1,1,1,0.0,44.11,0.0,74.7,1,0,96075
4902,0,0,0,0,24,1,0,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),56.35,1381.2,0,45,4,30.18,5128,0,Platina,0,0,DSL,40.367964,-122.937379,0,56.35,0,0,None,215,1,0,0,0,24,0,0.0,724.3199999999998,0.0,1381.2,0,1,96076
4903,0,0,0,0,5,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,90.8,455.5,1,25,56,1.49,5090,1,Red Bluff,0,0,Fiber Optic,40.186772,-122.388361,0,94.432,0,0,Offer E,26438,0,0,0,1,5,5,0.0,7.45,0.0,455.5,1,1,96080
4904,0,0,0,0,33,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,107.55,3645.5,0,39,12,49.69,4800,0,Round Mountain,1,0,DSL,40.923558,-122.059933,0,107.55,0,0,None,459,0,0,0,1,33,0,437.0,1639.77,0.0,3645.5,0,0,96084
4905,0,0,1,1,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.85,1158.85,0,48,0,11.81,6440,0,Scott Bar,0,0,NA,41.737961999999996,-123.07557,1,19.85,3,9,Offer B,88,0,0,1,0,58,0,0.0,684.98,0.0,1158.85,0,0,96085
4906,0,0,1,1,72,1,1,Fiber optic,1,1,1,0,Two year,1,Bank transfer (automatic),95.9,6954.15,0,26,59,11.85,4213,0,Seiad Valley,0,0,Fiber Optic,41.924174,-123.26078799999999,1,95.9,3,9,None,332,0,0,1,0,72,0,0.0,853.1999999999998,0.0,6954.15,1,1,96086
4907,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,23.85,1672.1,0,55,0,21.19,6166,0,Shasta,0,0,NA,40.617614,-122.51286100000002,1,23.85,0,4,None,528,0,0,1,0,71,0,0.0,1504.49,0.0,1672.1,0,0,96087
4908,0,1,0,0,28,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,106.15,3152.5,1,75,31,9.67,5030,1,Shingletown,1,0,DSL,40.497440999999995,-121.827524,0,110.39600000000002,0,0,Offer C,4231,0,0,0,0,28,2,977.0,270.76,0.0,3152.5,0,0,96088
4909,1,0,1,0,51,1,0,DSL,1,1,1,1,Two year,1,Credit card (automatic),83.85,4307.1,0,20,41,6.89,5703,0,Tehama,1,1,Fiber Optic,40.021786999999996,-122.127576,1,83.85,0,5,Offer B,405,1,0,1,1,51,0,176.59,351.39,0.0,4307.1,1,1,96090
4910,0,0,0,0,30,1,0,DSL,1,1,1,1,One year,0,Bank transfer (automatic),85.35,2530.4,1,59,4,43.01,2313,1,Trinity Center,1,0,Fiber Optic,41.081846999999996,-122.70054499999999,0,88.764,0,0,None,734,1,0,0,1,30,4,101.0,1290.3,0.0,2530.4,0,0,96091
4911,1,1,1,0,72,1,0,Fiber optic,1,1,0,0,Two year,1,Credit card (automatic),84.8,6141.65,0,77,2,5.51,4240,0,Vina,0,1,Cable,39.955164,-122.01856699999999,1,84.8,0,7,None,439,1,0,1,0,72,1,0.0,396.72,0.0,6141.65,0,1,96092
4912,1,1,0,0,36,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Electronic check,90.85,3186.7,1,69,25,23.33,5692,1,Weaverville,0,1,Cable,40.759401000000004,-122.93933700000001,0,94.484,0,0,Offer C,3749,0,2,0,0,36,3,797.0,839.8799999999999,0.0,3186.7,0,0,96093
4913,1,0,0,1,14,1,0,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),76.1,1054.8,0,24,52,36.73,2045,0,Weed,1,1,Cable,41.465121,-122.38094699999999,0,76.1,3,0,None,5896,1,0,0,1,14,1,548.0,514.2199999999998,0.0,1054.8,1,0,96094
4914,0,0,1,1,72,1,1,DSL,1,1,1,0,Two year,0,Mailed check,74.55,5430.65,0,61,30,21.84,4703,0,Whitmore,0,0,DSL,40.637105,-121.906949,1,74.55,3,9,None,843,1,0,1,0,72,1,0.0,1572.48,0.0,5430.65,0,1,96096
4915,0,0,1,1,22,0,No phone service,DSL,0,1,1,0,Month-to-month,0,Electronic check,39.2,849.9,0,53,19,0.0,3288,0,Yreka,0,0,Cable,41.764869,-122.67131599999999,1,39.2,1,4,None,9538,0,0,1,0,22,1,161.0,0.0,0.0,849.9,0,0,96097
4916,0,0,0,0,2,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,79.55,151.75,0,45,6,25.56,5965,0,Alturas,0,0,Fiber Optic,41.468877,-120.54229,0,79.55,0,0,Offer E,5096,0,2,0,0,2,2,0.0,51.12,0.0,151.75,0,1,96101
4917,0,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.6,299.4,0,48,0,39.87,3195,0,Blairsden Graeagle,0,0,NA,39.783747,-120.661032,0,19.6,0,0,None,1839,0,1,0,0,15,3,0.0,598.05,0.0,299.4,0,0,96103
4918,1,0,1,1,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.55,1086.75,0,40,0,28.96,5974,0,Cedarville,0,1,NA,41.505916,-120.152505,1,19.55,1,1,Offer B,857,0,0,1,0,51,0,0.0,1476.96,0.0,1086.75,0,0,96104
4919,1,0,1,0,70,0,No phone service,DSL,1,0,0,0,Two year,1,Credit card (automatic),39.15,2692.75,0,47,18,0.0,5840,0,Chilcoot,1,1,DSL,39.872961,-120.198876,1,39.15,0,1,None,650,1,0,1,0,70,0,48.47,0.0,0.0,2692.75,0,1,96105
4920,0,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.1,1389.6,0,45,0,31.03,5043,0,Clio,0,0,NA,39.745805,-120.580882,1,20.1,2,1,None,88,0,2,1,0,71,2,0.0,2203.13,0.0,1389.6,0,0,96106
4921,0,0,1,1,39,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),99.95,3767.4,0,35,53,24.38,4447,0,Coleville,0,0,Fiber Optic,38.42528,-119.47574099999999,1,99.95,3,1,None,1332,1,0,1,1,39,1,0.0,950.82,0.0,3767.4,0,1,96107
4922,0,0,1,1,61,1,1,DSL,1,1,0,0,Month-to-month,0,Electronic check,59.8,3641.5,0,27,30,26.7,5381,0,Davis Creek,0,0,Fiber Optic,41.750353999999994,-120.403885,1,59.8,1,1,Offer B,104,0,1,1,0,61,1,1092.0,1628.7,0.0,3641.5,1,0,96108
4923,0,0,0,0,52,1,0,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),49.75,2535.55,0,33,8,38.93,6334,0,Doyle,0,0,Fiber Optic,40.012675,-120.10185700000001,0,49.75,0,0,Offer B,1177,0,0,0,0,52,1,203.0,2024.36,0.0,2535.55,0,0,96109
4924,0,0,0,0,1,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,35.75,35.75,1,47,2,0.0,3351,1,Eagleville,0,0,Cable,41.280341,-120.15038100000001,0,37.18,0,0,Offer E,132,0,0,0,0,1,5,0.0,0.0,0.0,35.75,0,0,96110
4925,1,0,1,0,64,1,1,Fiber optic,1,0,1,1,One year,1,Mailed check,108.5,6880.85,0,27,71,4.01,4576,0,Fort Bidwell,1,1,Fiber Optic,41.932207,-120.13594099999999,1,108.5,0,1,Offer B,231,1,0,1,1,64,1,4885.0,256.64,0.0,6880.85,1,0,96112
4926,1,0,1,0,62,1,0,DSL,0,1,0,0,Two year,1,Credit card (automatic),60.15,3753.2,0,47,15,33.7,4404,0,Herlong,1,1,Fiber Optic,40.198234,-120.18088999999999,1,60.15,0,1,Offer B,946,1,0,1,0,62,1,0.0,2089.4,0.0,3753.2,0,1,96113
4927,1,0,1,0,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.05,637.55,0,64,0,11.38,2347,0,Janesville,0,1,NA,40.294034,-120.512622,1,19.05,0,1,None,3093,0,0,1,0,30,0,0.0,341.4000000000001,0.0,637.55,0,0,96114
4928,0,1,1,1,4,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,46.0,181.6,1,68,57,42.13,4797,1,Fallbrook,0,0,DSL,33.362575,-117.299644,1,47.84,3,1,Offer E,42239,0,0,1,0,4,6,104.0,168.52,0.0,181.6,0,0,92028
4929,1,1,1,0,63,1,0,DSL,1,1,1,1,One year,1,Bank transfer (automatic),84.0,5329.55,0,65,29,40.65,5688,0,Likely,1,1,Cable,41.266008,-120.49073100000001,1,84.0,0,1,None,277,1,0,1,1,63,2,154.56,2560.95,0.0,5329.55,0,1,96116
4930,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),44.55,44.55,0,27,82,23.04,5825,0,Litchfield,0,0,Fiber Optic,40.507272,-120.338228,0,44.55,0,0,Offer E,385,0,0,0,0,1,0,0.0,23.04,0.0,44.55,1,1,96117
4931,1,0,1,0,15,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,103.45,1539.8,0,59,13,18.6,5640,0,Loyalton,1,1,Fiber Optic,39.637471000000005,-120.22633799999998,1,103.45,0,1,None,1822,1,0,1,1,15,0,0.0,279.0,0.0,1539.8,0,1,96118
4932,1,0,1,1,27,1,0,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),80.65,2209.75,0,47,53,15.71,5856,0,Madeline,0,1,Fiber Optic,41.042003,-120.50608600000001,1,80.65,3,1,None,85,0,0,1,0,27,2,0.0,424.17,0.0,2209.75,0,1,96119
4933,0,0,0,1,4,0,No phone service,DSL,1,1,1,1,Month-to-month,1,Mailed check,57.2,223.75,0,31,52,0.0,2421,0,Markleeville,1,0,Fiber Optic,38.735789000000004,-119.85798,0,57.2,3,0,Offer E,957,0,0,0,1,4,0,116.0,0.0,0.0,223.75,0,0,96120
4934,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,110.75,7751.7,0,48,5,39.74,4848,0,Milford,1,0,Cable,40.181278999999996,-120.392967,1,110.75,0,1,None,481,0,0,1,1,72,1,0.0,2861.28,0.0,7751.7,0,1,96121
4935,1,1,1,0,45,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),24.7,1174.35,0,79,0,44.91,5644,0,Portola,0,1,NA,39.786755,-120.445626,1,24.7,0,5,None,4236,0,0,1,0,45,1,0.0,2020.95,0.0,1174.35,0,0,96122
4936,0,1,0,0,45,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,97.05,4385.05,0,71,4,12.67,4735,0,Ravendale,0,0,Cable,40.845738,-120.32221899999999,0,97.05,0,0,None,61,1,0,0,0,45,0,175.0,570.15,0.0,4385.05,0,0,96123
4937,0,0,0,0,36,1,0,DSL,1,1,1,0,One year,1,Mailed check,76.35,2606.35,0,33,8,44.87,4771,0,Calpine,1,0,Fiber Optic,39.672813,-120.456699,0,76.35,0,0,None,322,1,1,0,0,36,1,0.0,1615.32,0.0,2606.35,0,1,96124
4938,1,0,1,1,17,1,0,Fiber optic,1,0,1,0,Month-to-month,1,Electronic check,89.4,1539.45,1,54,24,19.19,2544,1,Sierra City,1,1,Fiber Optic,39.600599,-120.636358,1,92.976,0,1,None,348,0,0,1,0,17,0,369.0,326.23,0.0,1539.45,0,0,96125
4939,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,18.9,18.9,0,24,0,49.51,4480,0,Sierraville,0,1,NA,39.559709000000005,-120.34563899999999,0,18.9,0,0,Offer E,227,0,0,0,0,1,1,0.0,49.51,0.0,18.9,1,0,96126
4940,1,1,0,0,16,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.45,1261.35,0,70,5,22.02,5111,0,Standish,0,1,Fiber Optic,40.346634,-120.386422,0,74.45,0,0,Offer D,408,0,0,0,0,16,0,0.0,352.32,0.0,1261.35,0,1,96128
4941,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.8,58.15,1,33,0,15.12,4323,1,Susanville,0,1,NA,40.559177000000005,-120.612113,0,19.8,0,0,Offer E,19440,0,1,0,0,3,3,0.0,45.36,0.0,58.15,0,0,96130
4942,1,0,1,1,4,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.9,225.6,1,55,63,8.58,5691,1,Termo,0,1,Fiber Optic,41.027281,-120.669427,1,52.93600000000001,3,1,Offer E,72,0,1,1,0,4,2,142.0,34.32,0.0,225.6,0,0,96132
4943,0,0,1,0,71,1,0,DSL,1,1,1,1,Two year,1,Credit card (automatic),84.4,5969.3,0,33,26,3.09,5619,0,Topaz,1,0,Fiber Optic,38.636052,-119.48916200000001,1,84.4,0,0,None,116,1,0,0,1,71,0,1552.0,219.39,0.0,5969.3,0,0,96133
4944,1,0,1,1,10,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,24.4,253.9,0,27,0,4.16,4458,0,Tulelake,0,1,NA,41.813521,-121.49266599999999,1,24.4,1,4,None,2595,0,0,1,0,10,1,0.0,41.6,0.0,253.9,1,0,96134
4945,1,0,1,1,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.05,400,0,55,0,3.87,4328,0,Wendel,0,1,NA,40.345949,-120.08118700000001,1,20.05,1,4,None,162,0,0,1,0,20,1,0.0,77.4,0.0,400.0,0,0,96136
4946,1,0,0,0,4,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,81.0,340.85,1,25,65,21.62,3591,1,Westwood,0,1,Cable,40.271535,-121.01808700000001,0,84.24000000000002,0,0,Offer E,4158,0,0,0,1,4,1,222.0,86.48,0.0,340.85,1,0,96137
4947,1,0,0,0,26,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.35,2515.3,1,55,30,40.17,4997,1,Carnelian Bay,1,1,DSL,39.227434,-120.091806,0,102.284,0,0,None,1943,0,2,0,1,26,1,755.0,1044.42,0.0,2515.3,0,0,96140
4948,0,0,0,0,4,1,0,DSL,0,0,1,0,Month-to-month,0,Credit card (automatic),55.5,227.35,0,57,10,38.96,2328,0,Homewood,0,0,Cable,39.117018,-120.212535,0,55.5,0,0,Offer E,858,0,0,0,0,4,0,0.0,155.84,0.0,227.35,0,1,96141
4949,1,0,0,0,5,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Mailed check,51.0,305.95,1,20,65,0.0,4630,1,Tahoma,0,1,DSL,39.061227,-120.179546,0,53.04,0,0,None,1291,0,1,0,1,5,3,199.0,0.0,0.0,305.95,1,0,96142
4950,0,0,1,0,4,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,91.65,365.4,1,55,15,21.81,2140,1,Kings Beach,0,0,DSL,39.246654,-120.029273,1,95.316,0,1,Offer E,4806,0,1,1,0,4,3,55.0,87.24,0.0,365.4,0,0,96143
4951,1,1,1,0,29,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.3,2357.75,0,73,12,36.75,2217,0,Tahoe City,0,1,Cable,39.178337,-120.162806,1,84.3,0,7,Offer C,4002,0,0,1,1,29,0,0.0,1065.75,0.0,2357.75,0,1,96145
4952,1,0,0,0,2,1,0,Fiber optic,1,1,1,1,Month-to-month,0,Electronic check,100.2,198.5,0,49,15,22.56,4855,0,Olympic Valley,0,1,Fiber Optic,39.191796999999994,-120.212401,0,100.2,0,0,Offer E,942,0,0,0,1,2,2,0.0,45.12,0.0,198.5,0,1,96146
4953,0,0,0,0,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.4,554.25,0,30,0,15.06,2265,0,Tahoe Vista,0,0,NA,39.241240000000005,-120.05476499999999,0,19.4,0,0,None,678,0,0,0,0,29,1,0.0,436.74,0.0,554.25,0,0,96148
4954,1,0,0,1,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.85,90.85,1,47,7,1.13,5086,1,South Lake Tahoe,0,1,Fiber Optic,38.911577,-120.106169,0,94.484,0,0,Offer E,33038,0,0,0,1,1,4,0.0,1.13,0.0,90.85,0,0,96150
4955,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,69.4,69.4,1,62,22,38.53,2847,1,San Diego,0,1,DSL,32.957195,-117.202542,0,72.176,0,0,Offer E,28201,0,1,0,0,1,3,0.0,38.53,0.0,69.4,0,1,92130
4956,0,1,0,0,8,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),94.45,742.95,1,66,9,5.21,3676,1,Los Angeles,1,0,Cable,33.973616,-118.24902,0,98.228,0,0,Offer E,54492,0,1,0,0,8,3,0.0,41.68,0.0,742.95,0,1,90001
4957,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.4,251.65,0,56,0,46.92,2486,0,Los Angeles,0,1,NA,33.949255,-118.246978,0,20.4,0,0,None,44586,0,0,0,0,13,1,0.0,609.96,0.0,251.65,0,0,90002
4958,0,0,1,0,59,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,94.75,5597.65,0,60,14,16.39,5238,0,Los Angeles,0,0,Fiber Optic,33.964131,-118.272783,1,94.75,0,4,Offer B,58198,0,0,1,0,59,2,78.37,967.01,0.0,5597.65,0,1,90003
4959,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.15,20.15,1,55,0,3.09,4277,1,Los Angeles,0,0,NA,34.076259,-118.31071499999999,1,20.15,1,1,Offer E,67852,0,0,1,0,1,7,0.0,3.09,0.0,20.15,0,0,90004
4960,1,1,0,0,50,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.7,4816.7,1,65,12,18.92,4287,1,Los Angeles,0,1,Fiber Optic,34.059281,-118.30742,0,99.52799999999999,0,0,None,43019,0,1,0,1,50,4,0.0,946.0,0.0,4816.7,0,1,90005
4961,1,0,1,0,18,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),44.35,768.05,0,41,17,45.92,2935,0,Los Angeles,0,1,DSL,34.048013,-118.293953,1,44.35,0,10,Offer D,62784,0,0,1,0,18,0,131.0,826.5600000000002,0.0,768.05,0,0,90006
4962,0,0,1,1,17,1,0,DSL,1,1,1,1,Month-to-month,0,Mailed check,74.55,1215.8,0,22,47,44.9,4451,0,Los Angeles,0,0,Fiber Optic,34.027337,-118.28515,1,74.55,2,8,Offer D,45025,0,1,1,1,17,1,0.0,763.3,0.0,1215.8,1,1,90007
4963,1,0,1,0,47,1,0,DSL,0,1,1,1,Two year,0,Electronic check,73.6,3522.65,0,55,28,14.14,4795,0,Los Angeles,1,1,DSL,34.008293,-118.34676599999999,1,73.6,0,10,Offer B,30852,0,0,1,1,47,0,986.0,664.58,0.0,3522.65,0,0,90008
4964,0,0,0,0,26,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.95,1834.95,1,48,16,17.53,2934,1,Los Angeles,0,0,DSL,34.062125,-118.31570900000001,0,77.94800000000002,0,0,None,1957,0,0,0,0,26,3,294.0,455.78,0.0,1834.95,0,0,90010
4965,0,0,0,0,6,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,47.95,305.1,1,23,78,0.0,2240,1,Los Angeles,1,0,DSL,34.007090000000005,-118.25868100000001,0,49.868,0,0,Offer E,101215,0,1,0,1,6,4,238.0,0.0,0.0,305.1,1,0,90011
4966,1,0,1,1,19,1,1,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),50.1,910.45,0,51,13,9.47,5749,0,Los Angeles,0,1,DSL,34.065875,-118.23872800000001,1,50.1,2,10,Offer D,30596,0,0,1,0,19,3,118.0,179.93,0.0,910.45,0,0,90012
4967,0,0,0,0,3,1,1,DSL,0,0,1,0,Month-to-month,1,Electronic check,63.6,155.65,1,57,28,3.64,3155,1,Los Angeles,0,0,Cable,34.044639000000004,-118.24041299999999,0,66.14399999999999,0,0,Offer E,9732,1,1,0,0,3,2,44.0,10.92,0.0,155.65,0,0,90013
4968,0,1,1,1,68,0,No phone service,DSL,0,1,1,1,Two year,1,Electronic check,53.0,3656.25,0,65,23,0.0,5583,0,Los Angeles,1,0,Fiber Optic,34.043144,-118.251977,1,53.0,1,4,None,3524,0,0,1,1,68,0,84.09,0.0,0.0,3656.25,0,1,90014
4969,0,0,1,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.85,52,0,27,0,36.05,4107,0,Los Angeles,0,0,NA,34.039224,-118.26629299999999,1,19.85,0,8,Offer E,15140,0,0,1,0,2,2,0.0,72.1,0.0,52.0,1,0,90015
4970,1,0,0,0,7,0,No phone service,DSL,0,0,0,0,One year,1,Credit card (automatic),24.35,150.85,0,23,48,0.0,4665,0,Los Angeles,0,1,DSL,34.028331,-118.35433799999998,0,24.35,0,0,Offer E,46984,0,0,0,0,7,2,0.0,0.0,0.0,150.85,1,1,90016
4971,0,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.55,389.25,0,49,0,10.67,2386,0,Los Angeles,0,0,NA,34.052842,-118.264495,0,19.55,0,0,Offer D,20692,0,0,0,0,18,0,0.0,192.06,0.0,389.25,0,0,90017
4972,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.05,1873.7,0,46,0,44.84,6334,0,Los Angeles,0,0,NA,34.028735,-118.31723600000001,1,25.05,0,0,None,47143,0,0,0,0,71,1,0.0,3183.640000000001,0.0,1873.7,0,0,90018
4973,1,1,1,0,13,1,1,Fiber optic,1,1,0,1,Month-to-month,0,Credit card (automatic),93.8,1261,0,79,6,48.15,5870,0,Los Angeles,0,1,DSL,34.049841,-118.33846000000001,1,93.8,0,8,Offer D,67520,0,0,1,1,13,1,0.0,625.9499999999998,0.0,1261.0,0,1,90019
4974,1,0,0,0,3,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Mailed check,36.85,108.7,1,44,23,0.0,5825,1,San Diego,0,1,Fiber Optic,32.898613,-117.202937,0,38.32400000000001,0,0,Offer E,4258,1,1,0,0,3,1,25.0,0.0,0.0,108.7,0,0,92121
4975,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),103.75,7346.2,0,38,22,16.5,4655,0,Los Angeles,1,1,DSL,34.029043,-118.23950400000001,1,103.75,0,8,None,3012,0,0,1,1,72,0,1616.0,1188.0,0.0,7346.2,0,0,90021
4976,1,0,1,1,66,0,No phone service,DSL,0,1,1,1,Two year,1,Credit card (automatic),56.75,3708.4,0,35,25,0.0,5748,0,Los Angeles,1,1,Fiber Optic,34.02381,-118.156582,1,56.75,3,4,None,68701,0,0,1,1,66,2,927.0,0.0,0.0,3708.4,0,0,90022
4977,1,0,1,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.8,469.65,0,19,0,25.84,4654,0,Los Angeles,0,1,NA,34.017697,-118.200577,1,20.8,2,6,Offer C,47487,0,0,1,0,24,0,0.0,620.16,0.0,469.65,1,0,90023
4978,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.1,44.1,1,31,33,4.41,5955,1,Los Angeles,0,0,Fiber Optic,34.066303000000005,-118.435479,0,45.864,0,0,Offer E,44150,0,1,0,0,1,3,0.0,4.41,0.0,44.1,0,0,90024
4979,0,0,1,1,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.45,1385.85,0,20,0,31.53,5577,0,Los Angeles,0,0,NA,34.046174,-118.44633300000001,1,24.45,2,2,Offer B,41175,0,0,1,0,56,0,0.0,1765.68,0.0,1385.85,1,0,90025
4980,0,1,1,0,22,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),25.6,548.8,0,69,0,15.27,2628,0,Los Angeles,0,0,NA,34.078990999999995,-118.26380400000001,1,25.6,0,5,Offer D,73686,0,0,1,0,22,0,0.0,335.94,0.0,548.8,0,0,90026
4981,1,0,0,0,14,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,50.75,712.75,1,38,7,0.0,4883,1,Los Angeles,1,1,DSL,34.127194,-118.295647,0,52.78,0,0,Offer D,48727,0,2,0,1,14,3,50.0,0.0,0.0,712.75,0,0,90027
4982,0,1,1,0,61,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),104.4,6405,1,77,19,35.11,4412,1,Los Angeles,1,0,Cable,34.099869,-118.326843,1,108.576,0,1,None,30568,0,2,1,0,61,4,1217.0,2141.71,0.0,6405.0,0,0,90028
4983,0,1,1,0,40,0,No phone service,DSL,0,1,1,0,Month-to-month,1,Electronic check,39.3,1637.4,1,66,3,0.0,2296,1,Los Angeles,0,0,DSL,34.089953,-118.294824,1,40.872,0,1,None,41713,0,0,1,0,40,1,49.0,0.0,0.0,1637.4,0,0,90029
4984,0,0,0,0,42,1,0,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),59.65,2536.55,0,27,26,22.08,3048,0,Los Angeles,1,0,Fiber Optic,34.085807,-118.206617,0,59.65,0,0,Offer B,38415,0,0,0,0,42,0,660.0,927.36,0.0,2536.55,1,0,90031
4985,0,0,1,1,72,1,1,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),83.3,6042.7,0,28,69,24.48,4505,0,Los Angeles,1,0,Fiber Optic,34.078821000000005,-118.177576,1,83.3,3,3,None,46960,1,0,1,1,72,2,4169.0,1762.56,0.0,6042.7,1,0,90032
4986,0,0,0,0,12,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),79.55,958.25,0,47,16,21.93,3445,0,Los Angeles,0,0,Fiber Optic,34.050197999999995,-118.21094599999999,0,79.55,0,0,Offer D,49431,1,0,0,0,12,2,153.0,263.16,0.0,958.25,0,0,90033
4987,1,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.45,1730.65,0,24,0,33.61,4766,0,Los Angeles,0,1,NA,34.030578000000006,-118.39961299999999,1,24.45,0,2,None,58218,0,0,1,0,71,0,0.0,2386.31,0.0,1730.65,1,0,90034
4988,0,0,1,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.2,459.6,0,42,0,1.75,3656,0,Los Angeles,0,0,NA,34.051809000000006,-118.383843,1,19.2,0,10,Offer C,27799,0,0,1,0,26,0,0.0,45.5,0.0,459.6,0,0,90035
4989,0,0,0,1,7,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,29.8,201.95,0,33,19,0.0,4236,0,Los Angeles,0,0,DSL,34.070291,-118.34919099999999,0,29.8,2,0,None,32901,0,0,0,0,7,1,38.0,0.0,0.0,201.95,0,0,90036
4990,0,0,1,1,6,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.5,285.2,0,41,29,29.41,5450,0,Los Angeles,0,0,Fiber Optic,34.002642,-118.287596,1,45.5,1,1,None,56709,0,0,1,0,6,1,83.0,176.46,0.0,285.2,0,0,90037
4991,0,0,0,0,58,1,0,Fiber optic,1,1,1,1,One year,1,Electronic check,106.45,6145.85,1,57,13,14.99,5902,1,Los Angeles,1,0,Fiber Optic,34.088017,-118.327168,0,110.708,0,0,Offer B,32562,0,0,0,1,58,4,799.0,869.42,0.0,6145.85,0,0,90038
4992,1,0,1,0,51,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),30.05,1529.45,0,61,6,0.0,5045,0,Los Angeles,0,1,DSL,34.110845,-118.25959499999999,1,30.05,0,9,None,29310,0,0,1,0,51,0,92.0,0.0,0.0,1529.45,0,0,90039
4993,1,0,1,1,72,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),65.65,4664.5,0,32,16,0.0,4934,0,Los Angeles,1,1,DSL,33.994524,-118.149953,1,65.65,1,1,None,9805,1,0,1,1,72,0,0.0,0.0,0.0,4664.5,0,1,90040
4994,0,0,0,0,18,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,96.05,1740.7,1,23,29,35.7,5581,1,Los Angeles,0,0,Cable,34.137412,-118.20760700000001,0,99.89200000000001,0,0,Offer D,27866,0,2,0,1,18,1,0.0,642.6,0.0,1740.7,1,1,90041
4995,0,0,0,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),75.1,552.95,1,35,25,18.99,5514,1,Los Angeles,0,0,Cable,34.11572,-118.19275400000001,0,78.104,0,0,Offer E,64672,0,0,0,0,7,1,138.0,132.92999999999998,0.0,552.95,0,0,90042
4996,0,0,0,0,47,1,1,DSL,1,1,0,1,Two year,0,Mailed check,74.05,3496.3,0,56,3,45.67,2831,0,Los Angeles,0,0,Fiber Optic,33.988543,-118.33408100000001,0,74.05,0,0,None,44764,1,0,0,1,47,1,105.0,2146.49,0.0,3496.3,0,0,90043
4997,1,1,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.7,93.7,1,72,22,41.43,4618,1,Los Angeles,0,1,Fiber Optic,33.952714,-118.292061,0,46.48800000000001,0,0,Offer E,87383,0,0,0,0,2,4,21.0,82.86,0.0,93.7,0,0,90044
4998,1,1,0,0,62,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),110.75,7053.35,0,66,8,47.8,5166,0,Los Angeles,1,1,Cable,33.954017,-118.402447,0,110.75,0,0,None,39334,1,0,0,1,62,0,564.0,2963.6,0.0,7053.35,0,0,90045
4999,0,0,1,1,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.7,301.55,0,44,0,7.14,5293,0,Los Angeles,0,0,NA,34.108455,-118.362081,1,19.7,2,10,Offer D,49839,0,0,1,0,16,2,0.0,114.24,0.0,301.55,0,0,90046
5000,1,0,0,0,6,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),49.5,312.7,0,60,22,26.76,5552,0,Los Angeles,0,1,DSL,33.958149,-118.30844099999999,0,49.5,0,0,None,47107,1,0,0,0,6,0,69.0,160.56,0.0,312.7,0,0,90047
5001,1,0,0,0,19,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),55.0,1046.5,1,55,25,4.3,4539,1,Los Angeles,1,1,Cable,34.072945000000004,-118.37267,0,57.2,0,0,Offer D,21739,1,0,0,0,19,0,262.0,81.7,0.0,1046.5,0,0,90048
5002,0,0,1,1,69,0,No phone service,DSL,1,0,0,1,Two year,1,Credit card (automatic),43.95,2960.1,0,19,59,0.0,4479,0,Los Angeles,1,0,Fiber Optic,34.091829,-118.491244,1,43.95,1,7,None,33523,0,1,1,1,69,2,1746.0,0.0,0.0,2960.1,1,0,90049
5003,1,0,1,1,11,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.35,834.2,1,35,21,9.14,5075,1,Los Angeles,0,1,Cable,33.987945,-118.370442,1,77.324,0,1,Offer D,8115,0,2,1,0,11,6,0.0,100.54,0.0,834.2,0,1,90056
5004,0,0,1,0,64,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,111.15,6953.4,0,41,21,8.6,5455,0,Los Angeles,1,0,Fiber Optic,34.061918,-118.27793899999999,1,111.15,0,4,None,44004,1,0,1,1,64,2,0.0,550.4,0.0,6953.4,0,1,90057
5005,0,0,1,0,39,1,0,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),104.7,4134.85,1,35,8,9.51,2371,1,Los Angeles,1,0,Cable,34.001616999999996,-118.222274,1,108.88799999999999,0,1,None,3642,1,0,1,1,39,3,331.0,370.89,0.0,4134.85,0,0,90058
5006,0,0,0,0,15,1,1,DSL,1,0,0,0,Month-to-month,1,Mailed check,55.7,899.8,1,60,9,40.66,4519,1,Los Angeles,0,0,Cable,33.927254,-118.249826,0,57.928,0,0,Offer D,38128,0,0,0,0,15,5,0.0,609.9,0.0,899.8,0,1,90059
5007,1,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.6,541.5,0,33,0,13.36,2305,0,Los Angeles,0,1,NA,33.921279999999996,-118.27418600000001,0,20.6,0,0,Offer C,24511,0,0,0,0,25,1,0.0,334.0,0.0,541.5,0,0,90061
5008,0,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.65,116.85,0,43,0,29.09,3945,0,Los Angeles,0,0,NA,34.003553000000004,-118.30893300000001,0,19.65,0,0,None,29299,0,1,0,0,6,1,0.0,174.54,0.0,116.85,0,0,90062
5009,1,0,1,0,66,1,1,Fiber optic,1,1,1,1,One year,0,Bank transfer (automatic),115.8,7942.15,0,28,41,43.77,5845,0,Los Angeles,1,1,Fiber Optic,34.044271,-118.18523700000001,1,115.8,0,9,None,55668,1,0,1,1,66,0,3256.0,2888.82,0.0,7942.15,1,0,90063
5010,0,0,0,0,61,1,1,DSL,0,1,1,1,Two year,0,Credit card (automatic),88.65,5321.25,0,60,22,19.58,4730,0,Los Angeles,1,0,DSL,34.037251,-118.423573,0,88.65,0,0,None,24505,1,1,0,1,61,1,0.0,1194.38,0.0,5321.25,0,1,90064
5011,0,1,1,0,43,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,94.5,4156.8,0,76,22,3.66,4745,0,Los Angeles,0,0,Fiber Optic,34.108833000000004,-118.22971499999998,1,94.5,0,4,None,47534,0,0,1,0,43,1,0.0,157.38,0.0,4156.8,0,1,90065
5012,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.1,223.6,0,25,0,8.82,5179,0,Los Angeles,0,0,NA,34.002028,-118.430656,0,20.1,0,0,Offer D,55204,0,0,0,0,12,1,0.0,105.84,0.0,223.6,1,0,90066
5013,1,1,0,0,23,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Bank transfer (automatic),34.65,768.45,0,78,2,0.0,2307,0,Los Angeles,0,1,Fiber Optic,34.057496,-118.413959,0,34.65,0,0,None,2527,0,0,0,1,23,1,0.0,0.0,0.0,768.45,0,1,90067
5014,1,1,1,0,71,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Bank transfer (automatic),52.3,3765.05,0,73,28,0.0,5491,0,Los Angeles,1,1,Fiber Optic,34.137411,-118.328915,1,52.3,0,10,None,21728,0,0,1,1,71,1,105.42,0.0,0.0,3765.05,0,1,90068
5015,0,0,0,0,34,1,1,DSL,0,0,1,0,Month-to-month,0,Mailed check,65.0,2157.5,0,32,27,45.28,5567,0,West Hollywood,0,0,Fiber Optic,34.093781,-118.38106100000002,0,65.0,0,0,Offer C,20408,1,0,0,0,34,0,0.0,1539.52,0.0,2157.5,0,1,90069
5016,0,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.85,108.05,1,57,0,6.17,3799,1,Los Angeles,0,0,NA,34.052917,-118.255178,0,19.85,0,0,None,21,0,1,0,0,5,3,0.0,30.85,0.0,108.05,0,0,90071
5017,0,0,1,0,41,0,No phone service,DSL,0,1,0,0,One year,0,Mailed check,35.45,1391.65,0,59,17,0.0,2954,0,Los Angeles,0,0,DSL,34.102084000000005,-118.451629,1,35.45,0,10,None,10470,1,0,1,0,41,0,0.0,0.0,0.0,1391.65,0,1,90077
5018,0,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.7,1379.8,0,53,0,48.04,5451,0,Bell,0,0,NA,33.970343,-118.17136799999999,1,19.7,1,9,None,105285,0,0,1,0,72,0,0.0,3458.88,0.0,1379.8,0,0,90201
5019,1,1,0,0,14,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.6,1273.3,0,65,10,37.62,3502,0,Beverly Hills,0,1,DSL,34.099891,-118.41433799999999,0,95.6,0,0,None,21397,0,0,0,1,14,2,127.0,526.68,0.0,1273.3,0,0,90210
5020,0,0,0,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.85,810.45,0,53,0,2.32,3523,0,Beverly Hills,0,0,NA,34.063947,-118.38300100000001,0,19.85,0,0,None,8321,0,0,0,0,41,0,0.0,95.12,0.0,810.45,0,0,90211
5021,0,0,1,1,23,1,1,Fiber optic,1,0,0,0,One year,0,Credit card (automatic),81.85,1810.85,0,51,30,5.7,5939,0,Beverly Hills,0,0,Cable,34.062095,-118.401508,1,81.85,3,3,Offer D,11355,0,0,1,0,23,1,54.33,131.1,0.0,1810.85,0,1,90212
5022,1,0,1,1,71,1,0,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),109.3,7782.85,0,36,57,28.47,5737,0,Compton,1,1,Fiber Optic,33.88151,-118.234451,1,109.3,3,4,None,47305,1,0,1,1,71,1,0.0,2021.37,0.0,7782.85,0,1,90220
5023,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,70.3,1,57,12,15.92,5963,1,Compton,0,0,DSL,33.885811,-118.20645900000001,0,73.112,0,0,Offer E,51387,0,1,0,0,1,1,0.0,15.92,0.0,70.3,0,0,90221
5024,1,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.4,1797.1,0,40,0,4.15,6011,0,Compton,0,1,NA,33.912246,-118.236773,1,25.4,0,8,None,29825,0,0,1,0,72,1,0.0,298.8,0.0,1797.1,0,0,90222
5025,1,0,1,1,6,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.8,377.85,0,48,20,38.5,2651,0,Culver City,0,1,Fiber Optic,33.993990999999994,-118.39703999999999,1,69.8,3,9,None,31963,0,0,1,0,6,0,76.0,231.0,0.0,377.85,0,0,90230
5026,1,0,1,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.0,445.3,0,64,0,24.22,2170,0,Culver City,0,1,NA,34.019323,-118.391902,1,20.0,1,2,Offer D,15195,0,0,1,0,23,1,0.0,557.06,0.0,445.3,0,0,90232
5027,1,1,1,0,10,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,85.55,851.75,1,77,30,6.01,3336,1,Downey,0,1,DSL,33.956228,-118.120993,1,88.97200000000001,0,0,Offer D,24908,0,0,0,0,10,1,25.55,60.1,0.0,851.75,0,1,90240
5028,0,0,0,0,72,1,0,Fiber optic,1,1,1,1,Two year,1,Electronic check,109.9,7624.2,0,19,73,41.91,5234,0,Downey,1,0,Fiber Optic,33.940884000000004,-118.128628,0,109.9,0,0,None,40152,1,0,0,1,72,1,5566.0,3017.5199999999995,0.0,7624.2,1,0,90241
5029,0,0,1,0,7,1,0,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),50.3,355.1,0,19,53,33.24,2547,0,Downey,0,0,Fiber Optic,33.921793,-118.140588,1,50.3,0,7,None,42459,0,0,1,0,7,0,18.82,232.68,0.0,355.1,1,1,90242
5030,1,0,0,1,6,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Mailed check,94.5,575.45,1,53,19,16.58,3469,1,El Segundo,1,1,Cable,33.917145,-118.401554,0,98.28,0,0,Offer E,16041,0,3,0,1,6,3,109.0,99.48,0.0,575.45,0,0,90245
5031,1,0,1,1,9,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.5,906.85,0,33,16,36.94,2757,0,Gardena,0,1,DSL,33.890853,-118.29796699999999,1,101.5,1,1,None,47758,1,0,1,1,9,0,145.0,332.46,0.0,906.85,0,0,90247
5032,0,0,0,0,12,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.15,1057.55,0,52,6,34.73,4041,0,Gardena,0,0,Cable,33.876482,-118.284077,0,89.15,0,0,Offer D,9960,0,0,0,1,12,0,63.0,416.76,0.0,1057.55,0,0,90248
5033,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.4,19.4,0,43,0,23.97,2742,0,Gardena,0,0,NA,33.90139,-118.315697,0,19.4,0,0,None,26442,0,0,0,0,1,0,0.0,23.97,0.0,19.4,0,0,90249
5034,0,1,1,1,48,0,No phone service,DSL,0,1,0,0,One year,0,Bank transfer (automatic),29.9,1388.75,0,75,19,0.0,2617,0,Hawthorne,0,0,DSL,33.914775,-118.348083,1,29.9,2,0,None,93315,0,0,0,0,48,2,0.0,0.0,0.0,1388.75,0,1,90250
5035,1,0,0,0,20,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,78.8,1641.3,0,45,24,45.39,2317,0,Hermosa Beach,0,1,DSL,33.865320000000004,-118.396336,0,78.8,0,0,Offer D,18693,0,0,0,0,20,2,39.39,907.8,0.0,1641.3,0,1,90254
5036,0,1,1,0,16,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),85.35,1375.15,1,66,30,9.93,5769,1,Huntington Park,0,0,Cable,33.97803,-118.217141,1,88.764,0,1,Offer D,78114,0,0,1,0,16,0,413.0,158.88,0.0,1375.15,0,0,90255
5037,0,0,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,79.65,152.7,1,56,23,29.04,5082,1,Lawndale,0,0,DSL,33.88856,-118.35181299999999,0,82.83600000000001,0,0,Offer E,33300,0,1,0,0,2,4,35.0,58.08,0.0,152.7,0,0,90260
5038,0,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.3,185.2,0,25,0,45.42,4190,0,Lynwood,0,0,NA,33.923573,-118.20066899999999,0,19.3,0,0,Offer D,69850,0,1,0,0,10,1,0.0,454.2000000000001,0.0,185.2,1,0,90262
5039,0,1,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.6,195.05,1,80,33,31.91,4322,1,Malibu,0,0,Cable,34.037037,-118.705803,0,82.78399999999998,0,0,Offer E,11,0,1,0,0,2,4,64.0,63.82,0.0,195.05,0,0,90263
5040,1,0,1,1,20,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Mailed check,96.8,1826.7,0,32,23,42.06,3222,0,Malibu,0,1,Fiber Optic,34.074571999999996,-118.831181,1,96.8,3,7,Offer D,19630,1,0,1,0,20,0,420.0,841.2,0.0,1826.7,0,0,90265
5041,1,0,1,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.65,417.5,0,27,0,46.47,4147,0,Manhattan Beach,0,1,NA,33.889632,-118.39737,1,20.65,0,8,Offer D,33758,0,1,1,0,20,2,0.0,929.4,0.0,417.5,1,0,90266
5042,1,0,1,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.8,344.5,0,33,0,13.13,4464,0,Maywood,0,1,NA,33.988572,-118.18656499999999,1,19.8,1,1,Offer D,28094,0,0,1,0,19,3,0.0,249.47000000000003,0.0,344.5,0,0,90270
5043,1,1,0,0,19,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Electronic check,90.6,1660,1,68,28,28.12,2373,1,Pacific Palisades,0,1,Cable,34.079449,-118.54830600000001,0,94.22399999999999,0,0,Offer D,22548,0,3,0,0,19,4,465.0,534.28,0.0,1660.0,0,0,90272
5044,1,0,1,0,22,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,104.6,2180.55,0,53,3,49.66,2429,0,Palos Verdes Peninsula,0,1,Cable,33.788208000000004,-118.404955,1,104.6,0,1,Offer D,24979,1,0,1,1,22,1,6.54,1092.52,0.0,2180.55,0,1,90274
5045,0,0,0,0,35,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),80.05,2835.9,0,63,6,13.14,3999,0,Rancho Palos Verdes,0,0,DSL,33.753146,-118.36745900000001,0,80.05,0,0,Offer C,41263,1,0,0,0,35,2,170.0,459.9,0.0,2835.9,0,0,90275
5046,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,45.15,45.15,0,43,10,42.34,4131,0,Redondo Beach,0,0,Cable,33.830453000000006,-118.384565,0,45.15,0,0,None,34191,0,0,0,0,1,1,0.0,42.34,0.0,45.15,0,1,90277
5047,1,0,0,0,39,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),73.15,2730.85,0,43,24,8.69,3271,0,Redondo Beach,0,1,Fiber Optic,33.873395,-118.37019,0,73.15,0,0,Offer C,37322,0,0,0,0,39,0,655.0,338.91,0.0,2730.85,0,0,90278
5048,0,1,1,0,54,1,0,Fiber optic,0,0,1,1,One year,1,Electronic check,99.1,5437.1,0,68,17,22.05,4118,0,South Gate,1,0,Fiber Optic,33.944624,-118.19261499999999,1,99.1,0,1,None,96267,1,0,1,1,54,2,0.0,1190.7,0.0,5437.1,0,1,90280
5049,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.2,20.2,1,48,0,43.52,3061,1,Topanga,0,0,NA,34.115192,-118.61017,0,20.2,0,0,None,5451,0,0,0,0,1,1,0.0,43.52,0.0,20.2,0,0,90290
5050,1,0,1,0,66,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),106.05,6981.35,1,30,57,23.51,5602,1,Venice,1,1,DSL,33.991782,-118.479229,1,110.292,0,0,None,31021,0,1,0,1,66,3,3979.0,1551.66,0.0,6981.35,0,0,90291
5051,1,0,0,0,56,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Mailed check,105.35,5794.45,0,31,24,37.99,5680,0,Marina Del Rey,0,1,Cable,33.977468,-118.445475,0,105.35,0,0,None,18058,1,0,0,1,56,3,1391.0,2127.44,0.0,5794.45,0,0,90292
5052,1,0,0,1,18,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),45.65,747.2,0,58,28,34.07,4403,0,Playa Del Rey,0,1,Cable,33.947305,-118.43984099999999,0,45.65,2,0,Offer D,11264,0,0,0,0,18,0,209.0,613.26,0.0,747.2,0,0,90293
5053,0,0,1,1,16,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),79.95,1267.95,0,30,69,49.85,3855,0,Inglewood,0,0,Fiber Optic,33.956445,-118.35863400000001,1,79.95,2,1,Offer D,37527,0,0,1,0,16,0,0.0,797.6,0.0,1267.95,0,1,90301
5054,0,0,0,0,68,1,0,DSL,1,0,0,0,One year,1,Credit card (automatic),54.45,3674.95,0,45,27,17.41,6309,0,Inglewood,1,0,Fiber Optic,33.975332,-118.35525200000001,0,54.45,0,0,Offer A,30779,0,0,0,0,68,2,0.0,1183.88,0.0,3674.95,0,1,90302
5055,0,1,1,0,53,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.1,1275.6,0,79,0,19.03,5295,0,Inglewood,0,0,NA,33.936291,-118.33263899999999,1,25.1,0,1,None,27778,0,1,1,0,53,2,0.0,1008.59,0.0,1275.6,0,0,90303
5056,0,0,1,1,72,1,1,DSL,1,0,1,1,Two year,0,Credit card (automatic),84.7,5893.9,0,46,19,24.9,6375,0,Inglewood,1,0,Fiber Optic,33.936827,-118.359824,1,84.7,1,1,Offer A,28680,1,0,1,1,72,0,0.0,1792.8,0.0,5893.9,0,1,90304
5057,1,0,0,0,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.85,724.65,0,52,11,7.32,5212,0,Inglewood,0,1,DSL,33.958134,-118.330905,0,75.85,0,0,Offer E,13779,0,0,0,0,9,0,0.0,65.88,0.0,724.65,0,1,90305
5058,0,0,0,0,30,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,48.8,1536.75,0,37,13,10.74,4864,0,Santa Monica,0,0,Cable,34.015481,-118.49323100000001,0,48.8,0,0,Offer C,5221,0,0,0,0,30,2,19.98,322.2,0.0,1536.75,0,1,90401
5059,0,0,0,0,36,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.15,3615.6,1,54,8,13.35,4188,1,Santa Monica,0,0,Fiber Optic,34.035849,-118.50350800000001,0,103.116,0,0,None,11509,0,3,0,1,36,3,0.0,480.6,0.0,3615.6,0,1,90402
5060,0,0,0,0,18,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,35.2,607.3,0,45,11,0.0,5381,0,Santa Monica,1,0,DSL,34.031529,-118.491156,0,35.2,0,0,Offer D,23559,1,0,0,0,18,0,67.0,0.0,0.0,607.3,0,0,90403
5061,0,1,1,1,55,1,1,DSL,1,0,1,0,One year,0,Electronic check,76.25,4154.55,0,66,19,34.57,4319,0,Santa Monica,1,0,DSL,34.026334000000006,-118.474222,1,76.25,1,1,None,19975,1,0,1,0,55,1,789.0,1901.35,0.0,4154.55,0,0,90404
5062,0,0,1,0,39,0,No phone service,DSL,1,0,1,1,Month-to-month,0,Electronic check,55.9,2184.35,1,50,14,0.0,5632,1,Santa Monica,1,0,DSL,34.005439,-118.477507,1,58.136,0,3,None,26099,0,0,1,1,39,4,306.0,0.0,0.0,2184.35,0,0,90405
5063,1,0,0,0,21,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,82.35,1852.85,1,25,53,12.76,2902,1,Torrance,0,1,Fiber Optic,33.833698999999996,-118.31438700000001,0,85.64399999999998,0,0,Offer D,40705,0,2,0,1,21,1,982.0,267.96,0.0,1852.85,1,0,90501
5064,1,0,0,0,2,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),40.4,77.15,1,34,9,0.0,3620,1,Torrance,1,1,DSL,33.833181,-118.29206200000002,0,42.016000000000005,0,0,Offer E,17058,1,0,0,0,2,3,7.0,0.0,0.0,77.15,0,0,90502
5065,1,1,0,0,33,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),24.9,847.8,0,73,0,3.15,5756,0,Torrance,0,1,NA,33.840399,-118.353714,0,24.9,0,0,Offer C,41979,0,1,0,0,33,1,0.0,103.95,0.0,847.8,0,0,90503
5066,1,0,1,0,44,0,No phone service,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),54.3,2390.45,0,63,18,0.0,3222,0,Torrance,1,1,Fiber Optic,33.867257,-118.330794,1,54.3,0,1,None,31678,0,0,1,1,44,0,0.0,0.0,0.0,2390.45,0,1,90504
5067,0,0,1,1,30,1,0,DSL,1,0,0,1,Month-to-month,0,Bank transfer (automatic),66.3,1923.5,0,47,17,16.48,4631,0,Torrance,0,0,DSL,33.807882,-118.34795700000001,1,66.3,2,1,Offer C,34873,1,0,1,1,30,0,0.0,494.4,0.0,1923.5,0,1,90505
5068,0,0,1,0,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.9,1493.2,0,44,0,14.91,4030,0,Whittier,0,0,NA,34.007353,-118.03368300000001,1,20.9,0,0,Offer A,32050,0,0,0,0,71,0,0.0,1058.61,0.0,1493.2,0,0,90601
5069,0,0,0,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.35,338.1,1,42,10,29.11,2220,1,Whittier,0,0,DSL,33.972119,-118.02018799999999,0,78.36399999999998,0,0,Offer E,26265,0,1,0,0,4,1,34.0,116.44,0.0,338.1,0,0,90602
5070,1,0,0,1,35,1,0,Fiber optic,0,0,1,0,One year,1,Electronic check,85.15,3030.6,1,37,18,25.51,5928,1,Whittier,1,1,Cable,33.945318,-117.992066,0,88.55600000000003,0,0,None,19109,0,1,0,0,35,1,0.0,892.85,0.0,3030.6,0,1,90603
5071,1,0,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),75.35,75.35,0,32,9,38.89,3514,0,Whittier,1,1,Fiber Optic,33.929704,-118.01208000000001,1,75.35,0,1,Offer E,37887,0,0,1,0,1,0,0.0,38.89,0.0,75.35,0,0,90604
5072,1,1,1,0,23,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.45,2184.85,0,80,14,45.21,5883,0,Whittier,1,1,DSL,33.960891,-118.03222199999999,1,104.45,0,1,None,38181,0,0,1,1,23,2,306.0,1039.83,0.0,2184.85,0,0,90605
5073,0,0,0,1,22,0,No phone service,DSL,0,0,1,1,One year,1,Credit card (automatic),49.45,1031.4,0,55,29,0.0,5941,0,Whittier,1,0,DSL,33.976678,-118.065875,0,49.45,2,0,None,32148,0,1,0,1,22,1,29.91,0.0,0.0,1031.4,0,1,90606
5074,0,0,0,1,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.45,921.3,0,25,0,45.64,4170,0,Buena Park,0,0,NA,33.845706,-118.012204,0,19.45,1,0,None,44442,0,2,0,0,49,1,0.0,2236.36,0.0,921.3,1,0,90620
5075,0,0,1,1,42,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,92.15,3875.4,0,33,53,17.75,5697,0,Buena Park,1,0,Fiber Optic,33.874224,-117.99336799999999,1,92.15,3,10,None,33528,0,0,1,1,42,2,2054.0,745.5,0.0,3875.4,0,0,90621
5076,0,0,1,1,33,1,0,Fiber optic,0,0,1,1,One year,1,Electronic check,93.8,3124.5,1,48,30,20.02,5080,1,La Palma,1,0,Cable,33.850504,-118.039892,1,97.552,0,5,None,15505,0,0,1,1,33,2,937.0,660.66,0.0,3124.5,0,0,90623
5077,0,0,1,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.85,144.15,0,38,0,35.26,3973,0,Cypress,0,0,NA,33.818477,-118.038307,1,19.85,1,2,Offer E,47344,0,0,1,0,7,1,0.0,246.82,0.0,144.15,0,0,90630
5078,0,0,1,1,67,1,1,Fiber optic,1,0,0,1,One year,1,Bank transfer (automatic),100.25,6689,0,52,30,3.04,5588,0,La Habra,1,0,Cable,33.940619,-117.9513,1,100.25,3,10,Offer A,67354,1,0,1,1,67,1,2007.0,203.68,0.0,6689.0,0,0,90631
5079,1,0,0,0,15,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,95.7,1451.1,0,24,47,9.97,4999,0,La Mirada,0,1,Fiber Optic,33.902045,-118.00896100000001,0,95.7,0,0,None,47568,1,0,0,1,15,0,0.0,149.55,0.0,1451.1,1,1,90638
5080,1,0,1,0,67,1,1,Fiber optic,0,1,0,1,Two year,1,Electronic check,93.15,6368.2,0,42,11,17.4,4001,0,Montebello,1,1,Fiber Optic,34.015217,-118.10996200000001,1,93.15,0,5,Offer A,62425,0,0,1,1,67,2,701.0,1165.8,0.0,6368.2,0,0,90640
5081,1,0,1,1,53,1,0,DSL,1,1,1,0,Two year,1,Mailed check,69.7,3729.6,0,61,16,31.69,4590,0,Norwalk,0,1,Fiber Optic,33.905963,-118.08263000000001,1,69.7,2,3,None,103214,1,0,1,0,53,0,0.0,1679.5700000000004,0.0,3729.6,0,1,90650
5082,1,0,1,1,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.8,350.1,0,38,0,18.0,3243,0,Pico Rivera,0,1,NA,33.989523999999996,-118.089299,1,19.8,1,10,None,63288,0,0,1,0,21,1,0.0,378.0,0.0,350.1,0,0,90660
5083,0,0,1,1,40,1,0,DSL,1,1,0,1,Month-to-month,1,Mailed check,71.35,2847.2,0,30,48,29.14,5807,0,Santa Fe Springs,0,0,Fiber Optic,33.933565,-118.062611,1,71.35,2,4,None,16271,1,0,1,1,40,1,1367.0,1165.6,0.0,2847.2,0,0,90670
5084,0,0,1,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.75,452.35,0,49,0,45.35,2258,0,Stanton,0,0,NA,33.801869,-117.99506799999999,1,20.75,2,8,None,29694,0,1,1,0,22,1,0.0,997.7,0.0,452.35,0,0,90680
5085,1,0,0,0,39,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,40.6,1494.5,0,25,26,0.0,4436,0,Artesia,0,1,Fiber Optic,33.867593,-118.08063700000001,0,40.6,0,0,Offer C,16398,1,2,0,1,39,1,0.0,0.0,0.0,1494.5,1,1,90701
5086,1,0,0,0,45,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,20.4,930.45,1,49,0,25.4,5398,1,Cerritos,0,1,NA,33.8681,-118.067402,0,20.4,0,0,Offer B,51556,0,0,0,0,45,3,0.0,1143.0,0.0,930.45,0,0,90703
5087,0,0,1,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,41.85,0,35,0,5.42,5761,0,Avalon,0,0,NA,33.391181,-118.421305,1,20.35,0,3,Offer E,3699,0,0,1,0,2,1,0.0,10.84,0.0,41.85,0,0,90704
5088,0,0,1,1,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.75,1272.05,0,43,0,12.26,4235,0,Bellflower,0,0,NA,33.887676,-118.12728899999999,1,19.75,2,3,None,72893,0,0,1,0,57,0,0.0,698.8199999999998,0.0,1272.05,0,0,90706
5089,1,0,1,1,8,1,0,DSL,0,0,1,0,Month-to-month,1,Electronic check,54.4,475.1,0,49,57,1.56,4854,0,Harbor City,0,1,Fiber Optic,33.798266,-118.30023700000001,1,54.4,3,10,Offer E,24660,0,1,1,0,8,1,271.0,12.48,0.0,475.1,0,0,90710
5090,1,1,1,0,7,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Credit card (automatic),94.7,673.1,1,78,19,9.7,3591,1,Lakewood,0,1,Fiber Optic,33.840524,-118.148403,1,98.488,0,0,None,30173,0,0,0,1,7,1,0.0,67.89999999999999,0.0,673.1,0,1,90712
5091,1,0,0,0,6,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),30.5,208.7,1,47,15,0.0,4667,1,Lakewood,0,1,DSL,33.847755,-118.112532,0,31.72,0,0,Offer E,27563,0,2,0,0,6,1,0.0,0.0,0.0,208.7,0,1,90713
5092,0,0,1,1,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.45,150.75,0,30,0,5.84,4484,0,Lakewood,0,0,NA,33.841027000000004,-118.078097,1,20.45,1,3,Offer E,20890,0,0,1,0,7,0,0.0,40.88,0.0,150.75,0,0,90715
5093,1,0,0,0,49,1,1,DSL,0,0,1,0,Two year,1,Bank transfer (automatic),66.15,3199,0,49,13,17.77,6138,0,Hawaiian Gardens,0,1,DSL,33.830431,-118.07407099999999,0,66.15,0,0,None,14852,1,0,0,0,49,0,416.0,870.73,0.0,3199.0,0,0,90716
5094,0,0,0,0,65,1,1,Fiber optic,1,1,0,0,One year,1,Electronic check,89.85,5844.65,0,47,7,38.33,6421,0,Lomita,0,0,DSL,33.794209,-118.31735400000001,0,89.85,0,0,None,21065,1,0,0,0,65,0,409.0,2491.45,0.0,5844.65,0,0,90717
5095,0,0,0,0,55,1,0,DSL,0,0,0,0,One year,0,Bank transfer (automatic),45.05,2462.6,0,48,5,33.6,4055,0,Los Alamitos,0,0,Cable,33.794990000000006,-118.065591,0,45.05,0,0,None,21343,0,0,0,0,55,0,0.0,1848.0,0.0,2462.6,0,1,90720
5096,1,0,1,1,71,1,1,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),86.85,6263.8,0,28,59,10.11,6452,0,Paramount,1,1,Fiber Optic,33.897121999999996,-118.164432,1,86.85,3,10,Offer A,55306,1,0,1,1,71,1,3696.0,717.81,0.0,6263.8,1,0,90723
5097,1,0,0,0,35,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Mailed check,96.75,3403.4,0,62,23,39.87,5154,0,San Pedro,1,1,DSL,33.736387,-118.28436299999998,0,96.75,0,0,Offer C,58639,1,0,0,0,35,2,783.0,1395.4499999999996,0.0,3403.4,0,0,90731
5098,1,1,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,77.0,237.75,1,74,22,48.34,3128,1,San Pedro,0,1,Cable,33.744119,-118.31448,0,80.08,0,0,None,21279,0,1,0,0,3,3,52.0,145.02,0.0,237.75,0,0,90732
5099,0,0,0,1,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.1,221.35,1,62,0,33.06,4500,1,Seal Beach,0,0,NA,33.75462,-118.071128,0,20.1,3,0,Offer D,24180,0,0,0,0,11,4,0.0,363.66,0.0,221.35,0,0,90740
5100,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.3,75.3,1,53,3,26.06,2176,1,Sunset Beach,1,0,Cable,33.719221000000005,-118.073596,0,78.312,0,0,Offer E,1107,0,1,0,0,1,4,0.0,26.06,0.0,75.3,0,0,90742
5101,1,0,0,0,17,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Bank transfer (automatic),106.65,1672.1,0,29,59,38.78,2754,0,Surfside,1,1,DSL,33.728273,-118.08530400000001,0,106.65,0,0,None,174,1,0,0,0,17,1,98.65,659.26,0.0,1672.1,1,1,90743
5102,0,0,1,0,72,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),110.15,7881.2,0,20,85,23.7,4498,0,Wilmington,1,0,DSL,33.782068,-118.26226299999999,1,110.15,0,5,Offer A,53323,1,0,1,1,72,0,0.0,1706.4,0.0,7881.2,1,1,90744
5103,0,0,1,1,28,1,0,Fiber optic,1,0,0,1,One year,1,Bank transfer (automatic),82.85,2320.8,0,30,69,16.13,5802,0,Carson,0,0,Fiber Optic,33.822295000000004,-118.26411,1,82.85,1,4,Offer C,55486,0,0,1,1,28,0,0.0,451.64,0.0,2320.8,0,1,90745
5104,0,0,1,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.1,370.5,0,59,0,25.54,4329,0,Carson,0,0,NA,33.859171,-118.25227199999999,1,20.1,0,4,None,25566,0,0,1,0,18,1,0.0,459.72,0.0,370.5,0,0,90746
5105,0,1,1,0,40,1,0,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),99.2,4062.2,1,74,24,19.76,5098,1,Long Beach,0,0,Fiber Optic,33.752524,-118.21073700000001,1,103.16799999999999,0,1,None,38427,1,1,1,1,40,3,97.49,790.4000000000002,0.0,4062.2,0,1,90802
5106,0,0,0,0,52,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,59.45,3043.7,0,30,59,9.37,6107,0,Long Beach,1,0,Cable,33.760458,-118.129725,0,59.45,0,0,None,31352,0,0,0,1,52,2,1796.0,487.24,0.0,3043.7,0,0,90803
5107,0,0,1,0,47,1,0,DSL,0,1,1,0,Month-to-month,1,Bank transfer (automatic),58.6,2723.4,0,53,18,3.2,2613,0,Long Beach,0,0,Fiber Optic,33.783046999999996,-118.1486,1,58.6,0,8,None,43467,0,0,1,0,47,0,49.02,150.4,0.0,2723.4,0,1,90804
5108,0,0,0,0,23,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),49.7,1081.25,0,44,2,42.26,4790,0,Long Beach,1,0,Fiber Optic,33.864622,-118.179626,0,49.7,0,0,None,91664,0,0,0,0,23,0,0.0,971.98,0.0,1081.25,0,1,90805
5109,1,0,1,1,66,1,0,DSL,1,1,0,0,Two year,0,Mailed check,65.85,4097.05,0,59,30,26.91,5500,0,Long Beach,1,1,Cable,33.802664,-118.179971,1,65.85,2,10,Offer A,49647,1,0,1,0,66,1,0.0,1776.06,0.0,4097.05,0,1,90806
5110,0,0,0,0,8,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.5,632.2,0,22,41,17.3,5777,0,Long Beach,0,0,Fiber Optic,33.830099,-118.182239,0,73.5,0,0,None,31556,0,0,0,0,8,0,0.0,138.4,0.0,632.2,1,1,90807
5111,1,1,0,0,47,1,0,Fiber optic,1,0,0,1,Month-to-month,0,Mailed check,85.5,4042.3,1,65,22,36.58,3645,1,Long Beach,0,1,DSL,33.823943,-118.11133500000001,0,88.92,0,0,None,37417,0,1,0,1,47,3,889.0,1719.26,0.0,4042.3,0,0,90808
5112,0,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,164.85,1,62,0,48.22,5595,1,Long Beach,0,0,NA,33.819814,-118.222416,0,20.05,0,0,Offer E,35656,0,0,0,0,7,5,0.0,337.54,0.0,164.85,0,0,90810
5113,0,0,1,1,71,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),113.65,8166.8,0,23,41,4.32,6208,0,Long Beach,1,0,Fiber Optic,33.781086,-118.199049,1,113.65,2,2,Offer A,63136,1,0,1,1,71,2,0.0,306.72,0.0,8166.8,1,1,90813
5114,0,1,0,0,50,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,83.4,4113.7,0,65,22,47.99,4977,0,Long Beach,0,0,Cable,33.771612,-118.14386599999999,0,83.4,0,0,None,19034,0,0,0,0,50,2,905.0,2399.5,0.0,4113.7,0,0,90814
5115,1,0,1,0,46,1,0,DSL,1,1,0,0,Two year,0,Mailed check,65.65,3047.15,0,23,41,46.71,2680,0,Long Beach,1,1,DSL,33.797638,-118.11662,1,65.65,0,3,None,38902,1,0,1,0,46,2,1249.0,2148.66,0.0,3047.15,1,0,90815
5116,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.4,70.4,1,40,16,29.63,4238,1,Long Beach,0,1,DSL,33.778436,-118.118648,0,73.21600000000002,0,0,Offer E,425,0,1,0,0,1,1,0.0,29.63,0.0,70.4,0,1,90822
5117,0,0,0,0,66,0,No phone service,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),61.35,4193.4,0,25,73,0.0,4824,0,Altadena,1,0,DSL,34.196837,-118.14223600000001,0,61.35,0,0,Offer A,36243,1,0,0,1,66,1,3061.0,0.0,0.0,4193.4,1,0,91001
5118,0,0,1,0,42,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),85.9,3729.75,0,60,13,20.58,2219,0,Arcadia,1,0,Fiber Optic,34.137319,-118.02983700000001,1,85.9,0,8,None,30028,1,0,1,0,42,4,485.0,864.3599999999999,0.0,3729.75,0,0,91006
5119,0,0,0,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,75.65,399.45,0,62,6,29.75,2296,0,Arcadia,0,0,DSL,34.128284,-118.04773200000001,0,75.65,0,0,None,30933,1,0,0,0,5,0,0.0,148.75,0.0,399.45,0,1,91007
5120,1,0,1,1,7,1,0,DSL,1,0,0,0,One year,1,Electronic check,49.75,331.3,1,24,94,36.14,5651,1,Duarte,0,1,Fiber Optic,34.145695,-117.95982,1,51.74,0,4,Offer E,27414,0,1,1,1,7,2,311.0,252.98,0.0,331.3,1,0,91010
5121,1,0,0,0,29,1,1,DSL,0,1,0,1,One year,0,Credit card (automatic),70.9,1964.6,0,25,47,28.83,2064,0,La Canada Flintridge,1,1,Cable,34.234912,-118.153729,0,70.9,0,0,Offer C,20200,0,0,0,1,29,3,0.0,836.0699999999998,0.0,1964.6,1,1,91011
5122,0,0,1,1,27,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,49.85,1336.15,0,37,30,19.32,5580,0,Monrovia,0,0,DSL,34.1528,-118.000482,1,49.85,5,5,Offer C,41067,0,0,1,0,27,0,0.0,521.64,0.0,1336.15,0,1,91016
5123,0,1,0,0,15,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),75.3,1147.45,1,70,30,7.99,4526,1,Montrose,0,0,Fiber Optic,34.2112,-118.230625,0,78.312,0,0,None,7527,0,0,0,0,15,2,0.0,119.85,0.0,1147.45,0,1,91020
5124,0,0,1,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.1,486.05,0,25,0,4.57,5306,0,Sierra Madre,0,0,NA,34.168686,-118.057505,1,20.1,3,1,Offer C,10558,0,0,1,0,25,1,0.0,114.25,0.0,486.05,1,0,91024
5125,0,0,1,0,11,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.0,1078.9,1,64,20,25.67,2120,1,South Pasadena,0,0,DSL,34.110444,-118.156957,1,97.76,0,1,Offer D,23984,0,0,1,1,11,3,0.0,282.37,0.0,1078.9,0,1,91030
5126,1,0,1,0,57,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,103.05,5925.75,0,36,13,31.79,5586,0,Sunland,1,1,Cable,34.282703999999995,-118.312929,1,103.05,0,4,None,18752,1,0,1,0,57,0,770.0,1812.03,0.0,5925.75,0,0,91040
5127,1,0,0,0,67,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),118.35,7804.15,1,53,30,22.66,6255,1,Tujunga,1,1,Fiber Optic,34.296574,-118.24483899999998,0,123.084,0,0,None,26753,1,1,0,1,67,1,0.0,1518.22,0.0,7804.15,0,1,91042
5128,0,1,1,0,47,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,99.7,4747.2,0,73,7,2.98,4787,0,Pasadena,1,0,Cable,34.146634999999996,-118.139225,1,99.7,0,3,None,16812,0,0,1,1,47,0,332.0,140.06,0.0,4747.2,0,0,91101
5129,0,0,0,0,13,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,81.9,1028.9,0,47,19,34.18,2054,0,Pasadena,0,0,Fiber Optic,34.167465,-118.165327,0,81.9,0,0,None,27891,0,0,0,0,13,0,0.0,444.34,0.0,1028.9,0,1,91103
5130,1,0,0,0,8,0,No phone service,DSL,1,0,0,0,Month-to-month,1,Electronic check,30.45,226.45,1,55,4,0.0,4549,1,Pasadena,0,1,Fiber Optic,34.165383,-118.123752,0,31.668000000000003,0,0,Offer E,38460,0,2,0,0,8,3,9.0,0.0,0.0,226.45,0,0,91104
5131,0,0,1,0,44,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.1,4364.1,1,19,65,11.24,5606,1,Pasadena,0,0,DSL,34.13946,-118.16664899999999,1,99.944,0,4,None,10253,0,1,1,1,44,4,0.0,494.56,0.0,4364.1,1,1,91105
5132,1,0,1,1,71,1,1,DSL,1,0,1,0,One year,1,Electronic check,66.2,4692.55,0,42,26,37.03,4756,0,Pasadena,0,1,Fiber Optic,34.139402000000004,-118.128658,1,66.2,3,0,Offer A,23742,0,0,0,0,71,0,1220.0,2629.13,0.0,4692.55,0,0,91106
5133,1,1,1,0,24,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.25,2433.9,1,70,12,49.76,2104,1,Pasadena,1,1,Cable,34.159007,-118.08735300000001,1,108.42,0,3,Offer C,32369,0,1,1,1,24,3,292.0,1194.24,0.0,2433.9,0,0,91107
5134,1,1,0,0,15,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.2,1217.25,1,75,6,12.08,4958,1,San Marino,0,1,Fiber Optic,34.122671000000004,-118.11291100000001,0,83.40799999999999,0,0,None,13158,0,0,0,0,15,5,0.0,181.2,0.0,1217.25,0,1,91108
5135,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.75,19.75,0,57,0,37.62,3666,0,Glendale,0,0,NA,34.17051,-118.28946299999998,0,19.75,0,0,None,23981,0,0,0,0,1,1,0.0,37.62,0.0,19.75,0,0,91201
5136,1,1,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,72.6,154.3,0,73,30,15.19,5098,0,Glendale,0,1,DSL,34.167926,-118.26753899999999,0,72.6,0,0,None,21990,0,0,0,0,2,0,0.0,30.38,0.0,154.3,0,1,91202
5137,1,1,0,0,55,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,116.5,6382.55,0,70,10,29.3,4222,0,Glendale,1,1,DSL,34.153338,-118.262974,0,116.5,0,0,None,14493,1,2,0,0,55,2,0.0,1611.5,0.0,6382.55,0,1,91203
5138,1,1,0,0,71,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,106.8,7623.2,0,67,21,34.8,6423,0,Glendale,0,1,Fiber Optic,34.136306,-118.26036,0,106.8,0,0,None,17015,1,1,0,0,71,1,0.0,2470.8,0.0,7623.2,0,1,91204
5139,1,0,1,1,50,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.95,1261.45,0,33,0,22.3,6019,0,Glendale,0,1,NA,34.13658,-118.24583899999999,1,24.95,1,3,None,41390,0,0,1,0,50,1,0.0,1115.0,0.0,1261.45,0,0,91205
5140,1,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.25,89.25,0,49,2,16.64,5579,0,Glendale,0,1,DSL,34.162515,-118.203869,0,89.25,0,0,None,31297,0,1,0,1,1,1,0.0,16.64,0.0,89.25,0,1,91206
5141,1,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.25,86.05,0,32,0,21.01,3056,0,Glendale,0,1,NA,34.182378,-118.262922,0,19.25,0,0,None,9864,0,0,0,0,5,2,0.0,105.05,0.0,86.05,0,0,91207
5142,0,0,0,0,66,1,1,Fiber optic,1,1,1,0,One year,1,Bank transfer (automatic),104.55,6779.05,0,44,26,16.39,4494,0,Glendale,1,0,DSL,34.195386,-118.23850800000001,0,104.55,0,0,Offer A,16910,1,0,0,0,66,0,1763.0,1081.74,0.0,6779.05,0,0,91208
5143,0,0,1,1,49,1,0,DSL,1,1,1,1,One year,1,Mailed check,87.2,4345,0,32,23,33.07,4567,0,La Crescenta,1,0,Fiber Optic,34.239636,-118.245259,1,87.2,2,4,None,29110,1,0,1,1,49,1,0.0,1620.43,0.0,4345.0,0,1,91214
5144,0,1,1,0,3,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,30.75,82.85,0,75,3,0.0,4133,0,Agoura Hills,0,0,Fiber Optic,34.129058,-118.75978799999999,1,30.75,0,7,None,25303,0,0,1,0,3,0,2.0,0.0,0.0,82.85,0,0,91301
5145,1,0,1,1,66,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),25.7,1714.55,0,32,0,42.84,5517,0,Calabasas,0,1,NA,34.130860999999996,-118.68346000000001,1,25.7,3,3,Offer A,23661,0,0,1,0,66,0,0.0,2827.44,0.0,1714.55,0,0,91302
5146,1,0,0,1,11,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,86.2,893.2,0,31,10,5.84,3157,0,Canoga Park,0,1,Fiber Optic,34.19829,-118.602203,0,86.2,2,0,None,23519,0,0,0,1,11,3,0.0,64.24,0.0,893.2,0,1,91303
5147,1,0,0,0,28,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),30.1,810.85,0,29,48,0.0,2653,0,Canoga Park,0,1,DSL,34.224377000000004,-118.63265600000001,0,30.1,0,0,Offer C,49242,1,0,0,0,28,2,0.0,0.0,0.0,810.85,1,1,91304
5148,1,0,1,0,65,1,1,Fiber optic,1,1,1,0,Two year,1,Electronic check,99.35,6347.55,0,31,20,30.44,6300,0,Winnetka,1,1,Cable,34.209532,-118.57756299999998,1,99.35,0,9,None,43857,0,0,1,0,65,1,0.0,1978.6,0.0,6347.55,0,1,91306
5149,0,0,0,0,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.2,1123.65,0,45,0,24.03,4937,0,West Hills,0,0,NA,34.199787,-118.68493000000001,0,19.2,0,0,None,23637,0,0,0,0,62,2,0.0,1489.86,0.0,1123.65,0,0,91307
5150,0,0,1,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.1,43.15,0,38,0,32.86,4158,0,Chatsworth,0,0,NA,34.294142,-118.60388300000001,1,20.1,0,9,None,35325,0,0,1,0,2,1,0.0,65.72,0.0,43.15,0,0,91311
5151,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.35,35.1,0,57,0,2.46,3746,0,Encino,0,0,NA,34.150354,-118.51829199999999,0,20.35,0,0,None,27614,0,0,0,0,2,0,0.0,4.92,0.0,35.1,0,0,91316
5152,0,0,1,1,55,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.65,1388,0,36,0,1.44,4466,0,Newbury Park,0,0,NA,34.172071,-118.946262,1,25.65,3,1,Offer B,37779,0,0,1,0,55,2,0.0,79.2,0.0,1388.0,0,0,91320
5153,1,1,1,0,41,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,94.55,3851.45,0,65,2,46.46,4914,0,Newhall,0,1,Fiber Optic,34.370378,-118.50411799999999,1,94.55,0,8,Offer B,30742,0,1,1,1,41,2,7.7,1904.86,0.0,3851.45,0,1,91321
5154,0,0,1,1,17,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,104.2,1743.5,1,38,16,4.91,2365,1,Northridge,1,0,Cable,34.238208,-118.55028999999999,1,108.368,0,1,Offer D,25751,0,0,1,1,17,1,279.0,83.47,0.0,1743.5,0,0,91324
5155,0,0,0,0,30,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),94.4,2638.1,0,64,27,2.67,4584,0,Northridge,0,0,Fiber Optic,34.236683,-118.51758799999999,0,94.4,0,0,None,32307,1,0,0,1,30,0,712.0,80.1,0.0,2638.1,0,0,91325
5156,1,0,0,0,17,1,0,DSL,1,1,0,0,One year,0,Mailed check,56.1,946.95,0,58,15,36.47,5025,0,Porter Ranch,0,1,Fiber Optic,34.281911,-118.55621799999999,0,56.1,0,0,None,28067,0,0,0,0,17,0,142.0,619.99,0.0,946.95,0,0,91326
5157,0,0,1,1,16,1,0,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),68.25,1114.85,0,32,30,20.12,3559,0,Pacoima,0,0,DSL,34.255441999999995,-118.421314,1,68.25,1,10,None,97318,1,0,1,1,16,0,33.45,321.92,0.0,1114.85,0,1,91331
5158,1,0,0,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.75,1777.6,0,25,0,29.29,5398,0,Reseda,0,1,NA,34.200175,-118.540958,0,24.75,0,0,Offer A,68018,0,0,0,0,72,1,0.0,2108.88,0.0,1777.6,1,0,91335
5159,1,0,0,0,9,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.25,684.85,0,48,3,34.75,2062,0,San Fernando,0,1,Fiber Optic,34.286131,-118.435969,0,76.25,0,0,None,33389,0,0,0,0,9,0,0.0,312.75,0.0,684.85,0,1,91340
5160,0,0,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,74.35,74.35,0,43,4,24.41,4237,0,Sylmar,0,0,DSL,34.321621,-118.399841,0,74.35,0,0,None,81986,0,0,0,0,1,0,0.0,24.41,0.0,74.35,0,1,91342
5161,1,0,0,1,23,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,54.15,1312.45,0,64,27,8.4,2496,0,North Hills,0,1,Fiber Optic,34.238802,-118.48229599999999,0,54.15,1,0,None,57017,1,1,0,0,23,1,0.0,193.2,0.0,1312.45,0,1,91343
5162,1,0,0,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.45,159.2,0,28,0,1.95,4119,0,Granada Hills,0,1,NA,34.291273,-118.505104,0,19.45,3,0,None,48867,0,0,0,0,8,2,0.0,15.6,0.0,159.2,1,0,91344
5163,1,0,1,1,19,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Mailed check,34.95,610.2,0,23,52,0.0,3422,0,Mission Hills,0,1,Fiber Optic,34.266389000000004,-118.459744,1,34.95,1,3,None,17112,0,0,1,0,19,0,0.0,0.0,0.0,610.2,1,1,91345
5164,0,0,0,0,7,1,1,DSL,1,0,0,0,Month-to-month,1,Electronic check,53.65,404.35,0,46,17,40.42,4389,0,Santa Clarita,0,0,Fiber Optic,34.502432,-118.41458999999999,0,53.65,0,0,Offer E,40077,0,0,0,0,7,1,69.0,282.94,0.0,404.35,0,0,91350
5165,1,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.65,69.65,1,70,2,7.23,5844,1,Canyon Country,0,1,Fiber Optic,34.422519,-118.420717,0,72.436,0,0,None,59259,0,0,0,0,1,5,0.0,7.23,0.0,69.65,0,0,91351
5166,1,0,0,0,61,1,1,Fiber optic,1,0,1,1,One year,0,Electronic check,104.0,6363.45,0,24,48,45.69,4344,0,Sun Valley,1,1,Cable,34.231053,-118.338307,0,104.0,0,0,Offer B,46639,0,0,0,1,61,1,305.45,2787.09,0.0,6363.45,1,1,91352
5167,0,0,1,0,57,1,0,DSL,1,1,1,0,Two year,1,Credit card (automatic),70.35,4124.65,0,32,24,48.0,5779,0,Valencia,0,0,Cable,34.457005,-118.57372600000001,1,70.35,0,1,Offer B,17846,1,0,1,0,57,2,0.0,2736.0,0.0,4124.65,0,1,91354
5168,1,0,0,0,9,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.8,713.1,1,39,8,20.34,3890,1,Valencia,0,1,Cable,34.43987,-118.644609,0,84.03200000000001,0,0,None,24977,0,0,0,1,9,2,57.0,183.06,0.0,713.1,0,0,91355
5169,1,0,0,1,15,1,0,DSL,1,0,0,1,One year,0,Mailed check,64.85,950.75,0,31,29,43.69,4442,0,Tarzana,1,1,DSL,34.157137,-118.548511,0,64.85,3,0,None,27424,0,0,0,1,15,1,276.0,655.3499999999998,0.0,950.75,0,0,91356
5170,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,19.65,0,42,0,23.67,4639,0,Thousand Oaks,0,0,NA,34.214054,-118.88108999999999,0,19.65,0,0,Offer E,42526,0,0,0,0,1,0,0.0,23.67,0.0,19.65,0,0,91360
5171,0,0,1,0,12,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),45.9,505.95,0,39,4,30.79,5790,0,Westlake Village,0,0,Fiber Optic,34.130992,-118.894673,1,45.9,0,0,None,18735,0,0,0,0,12,0,0.0,369.48,0.0,505.95,0,1,91361
5172,1,0,0,0,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.0,1149.65,0,48,0,27.3,6094,0,Thousand Oaks,0,1,NA,34.191842,-118.822796,0,20.0,0,0,Offer B,33057,0,0,0,0,54,2,0.0,1474.2,0.0,1149.65,0,0,91362
5173,1,0,1,1,4,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.8,169.65,0,40,19,25.9,2114,0,Woodland Hills,0,1,Cable,34.153733,-118.59340800000001,1,44.8,2,1,Offer E,25988,0,0,1,0,4,1,3.22,103.6,0.0,169.65,0,1,91364
5174,0,0,0,0,7,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,80.3,526.7,1,21,46,39.21,3949,1,Woodland Hills,0,0,DSL,34.178067999999996,-118.61571399999998,0,83.512,0,0,None,36123,0,0,0,1,7,3,242.0,274.47,0.0,526.7,1,0,91367
5175,0,0,1,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.35,393.15,0,23,0,27.96,4390,0,Oak Park,0,0,NA,34.19225,-118.77687399999999,1,20.35,0,1,None,14814,0,0,1,0,20,2,0.0,559.2,0.0,393.15,1,0,91377
5176,0,0,0,1,26,0,No phone service,DSL,1,0,0,1,Month-to-month,0,Mailed check,45.8,1147,0,51,19,0.0,3287,0,Stevenson Ranch,0,0,Cable,34.364153,-118.615583,0,45.8,2,0,None,9937,1,0,0,1,26,1,0.0,0.0,0.0,1147.0,0,1,91381
5177,1,1,1,0,36,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.1,3021.6,1,71,16,31.65,2987,1,Castaic,0,1,DSL,34.506627,-118.699048,1,87.464,0,1,Offer C,22177,0,0,1,0,36,2,483.0,1139.4,0.0,3021.6,0,0,91384
5178,0,0,1,0,53,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),108.95,5718.2,0,36,20,18.0,4163,0,Van Nuys,1,0,Fiber Optic,34.178483,-118.43179099999999,1,108.95,0,1,Offer B,40376,1,0,1,1,53,2,1144.0,954.0,0.0,5718.2,0,0,91401
5179,1,0,0,0,3,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,69.35,191.35,1,48,7,35.64,3520,1,Fallbrook,0,1,Cable,33.362575,-117.299644,0,72.124,0,0,None,42239,1,0,0,1,3,2,13.0,106.92,0.0,191.35,0,0,92028
5180,0,0,0,0,68,0,No phone service,DSL,1,1,1,1,Two year,0,Credit card (automatic),64.35,4539.6,0,38,28,0.0,4146,0,Sherman Oaks,1,0,DSL,34.147149,-118.463365,0,64.35,0,0,Offer A,22085,1,0,0,1,68,1,0.0,0.0,0.0,4539.6,0,1,91403
5181,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),90.8,6397.6,0,64,26,20.63,5028,0,Van Nuys,1,1,Fiber Optic,34.202494,-118.448048,1,90.8,2,1,Offer A,51348,1,0,1,1,72,1,1663.0,1485.36,0.0,6397.6,0,0,91405
5182,1,0,0,0,12,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),24.95,280.4,0,61,0,25.57,4443,0,Van Nuys,0,1,NA,34.195685,-118.490752,0,24.95,0,0,Offer D,50047,0,0,0,0,12,1,0.0,306.8400000000001,0.0,280.4,0,0,91406
5183,0,1,1,1,34,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,79.6,2718.3,1,79,16,25.84,3980,1,Van Nuys,0,0,Cable,34.178470000000004,-118.45947199999999,1,82.78399999999998,0,1,Offer C,23646,0,1,1,0,34,3,0.0,878.56,0.0,2718.3,0,1,91411
5184,0,0,1,0,68,1,1,Fiber optic,1,1,0,0,Two year,1,Bank transfer (automatic),84.7,5711.05,0,52,4,7.87,5520,0,Sherman Oaks,0,0,Fiber Optic,34.146957,-118.432138,1,84.7,0,1,Offer A,29387,0,0,1,0,68,0,0.0,535.16,0.0,5711.05,0,1,91423
5185,0,0,0,1,50,1,0,DSL,1,0,1,0,One year,1,Credit card (automatic),70.8,3478.15,0,25,71,37.52,4798,0,Encino,1,0,DSL,34.152875,-118.486056,0,70.8,2,0,Offer B,13129,1,0,0,0,50,3,0.0,1876.0,0.0,3478.15,1,1,91436
5186,0,1,0,0,1,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,36.45,36.45,1,79,29,0.0,5303,1,Burbank,0,0,Cable,34.188339,-118.30094199999999,0,37.908,0,0,None,18112,0,1,0,0,1,5,0.0,0.0,0.0,36.45,0,1,91501
5187,0,1,0,0,41,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.4,4133.95,0,78,15,6.33,4477,0,Burbank,1,0,Fiber Optic,34.177267,-118.31003,0,104.4,0,0,Offer B,11517,0,0,0,0,41,0,620.0,259.53000000000003,0.0,4133.95,0,0,91502
5188,1,1,1,0,30,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.5,2917.65,0,79,24,48.02,4828,0,Burbank,0,1,Fiber Optic,34.213049,-118.317651,1,101.5,0,1,Offer C,25882,1,0,1,0,30,1,0.0,1440.6,0.0,2917.65,0,1,91504
5189,1,0,0,0,1,1,1,DSL,0,1,0,0,Month-to-month,0,Electronic check,54.3,54.3,0,62,24,34.02,3259,0,Burbank,0,1,DSL,34.174215000000004,-118.345928,0,54.3,0,0,Offer E,29245,0,0,0,0,1,0,0.0,34.02,0.0,54.3,0,0,91505
5190,1,1,1,1,29,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,103.95,2964.8,0,69,19,49.36,3733,0,Burbank,1,1,Fiber Optic,34.169706,-118.323548,1,103.95,1,1,Offer C,18539,0,0,1,0,29,2,0.0,1431.44,0.0,2964.8,0,1,91506
5191,0,0,1,1,23,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),91.1,2198.3,0,20,51,27.97,5991,0,North Hollywood,1,0,Fiber Optic,34.1692,-118.372498,1,91.1,2,1,Offer D,36625,1,0,1,1,23,3,112.11,643.31,0.0,2198.3,1,1,91601
5192,1,0,0,1,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.95,1189.9,0,49,0,16.59,5316,0,North Hollywood,0,1,NA,34.15136,-118.36478600000001,0,19.95,2,0,Offer B,16996,0,0,0,0,60,2,0.0,995.4,0.0,1189.9,0,0,91602
5193,0,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),26.45,1914.5,0,21,0,22.22,5534,0,Studio City,0,0,NA,34.139082,-118.39275,1,26.45,0,1,Offer A,26157,0,0,1,0,72,0,0.0,1599.84,0.0,1914.5,1,0,91604
5194,1,0,0,1,22,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.4,2001.5,1,39,13,39.58,5438,1,North Hollywood,1,1,DSL,34.207295,-118.40002199999999,0,92.976,0,0,Offer D,57146,0,1,0,0,22,2,260.0,870.76,0.0,2001.5,0,0,91605
5195,1,0,0,0,72,1,0,DSL,1,1,1,0,Two year,1,Bank transfer (automatic),75.1,5336.35,0,32,22,15.03,6284,0,North Hollywood,1,1,DSL,34.187599,-118.387125,0,75.1,0,0,Offer A,45358,1,0,0,0,72,1,0.0,1082.16,0.0,5336.35,0,1,91606
5196,0,1,0,0,66,1,1,Fiber optic,0,1,1,1,One year,0,Bank transfer (automatic),108.1,7238.6,0,72,28,3.57,4722,0,Valley Village,1,0,Cable,34.165783000000005,-118.399795,0,108.1,0,0,None,27453,0,0,0,0,66,0,2027.0,235.62,0.0,7238.6,0,0,91607
5197,0,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,110.15,7998.8,0,54,24,12.85,5065,0,Rancho Cucamonga,1,0,Fiber Optic,34.132275,-117.611478,1,110.15,0,7,Offer A,39064,1,0,1,1,72,0,191.97,925.2,0.0,7998.8,0,1,91701
5198,0,1,1,0,47,1,1,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,80.35,3825.85,1,73,8,38.31,5915,1,Azusa,0,0,Cable,34.174493,-117.87068000000001,1,83.564,0,1,None,57775,0,1,1,0,47,2,306.0,1800.5700000000004,0.0,3825.85,0,0,91702
5199,0,0,0,0,51,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,111.5,5703.25,0,19,82,43.79,4363,0,Baldwin Park,1,0,Fiber Optic,34.098275,-117.967399,0,111.5,0,0,Offer B,76890,1,0,0,1,51,0,4677.0,2233.29,0.0,5703.25,1,0,91706
5200,0,0,1,1,70,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,106.5,7397,0,47,19,5.93,6319,0,Chino Hills,1,0,Cable,33.942895,-117.72564399999999,1,106.5,1,2,Offer A,66754,0,0,1,1,70,0,1405.0,415.1,0.0,7397.0,0,0,91709
5201,1,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,19.9,164.6,0,28,0,4.02,3643,0,Chino,0,1,NA,33.990646000000005,-117.663025,0,19.9,0,0,None,75319,0,0,0,0,9,2,0.0,36.17999999999999,0.0,164.6,1,0,91710
5202,1,0,1,1,59,1,1,Fiber optic,1,1,1,1,Two year,1,Mailed check,111.1,6555.2,0,40,57,46.1,4952,0,Claremont,0,1,DSL,34.127621000000005,-117.717863,1,111.1,3,1,Offer B,34716,1,0,1,1,59,0,0.0,2719.9,0.0,6555.2,0,1,91711
5203,1,0,0,1,3,1,0,DSL,0,0,1,1,Month-to-month,0,Mailed check,70.7,225.65,0,44,17,25.04,2584,0,Covina,0,1,DSL,34.097345000000004,-117.90673600000001,0,70.7,1,0,Offer E,33817,1,0,0,1,3,1,0.0,75.12,0.0,225.65,0,1,91722
5204,1,1,1,0,38,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.85,955.75,0,69,30,0.0,3511,0,Covina,0,1,Cable,34.084747,-117.886844,1,24.85,0,2,Offer C,17554,0,2,1,0,38,2,28.67,0.0,0.0,955.75,0,1,91723
5205,0,0,0,0,37,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Bank transfer (automatic),91.2,3382.3,0,52,30,11.73,5135,0,Covina,1,0,Fiber Optic,34.081109999999995,-117.853935,0,91.2,0,0,None,25068,0,0,0,0,37,2,1015.0,434.01,0.0,3382.3,0,0,91724
5206,1,0,0,0,37,1,0,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),65.6,2313.8,0,35,30,38.43,3183,0,Rancho Cucamonga,1,1,DSL,34.100970000000004,-117.57882,0,65.6,0,0,None,51970,1,0,0,0,37,1,694.0,1421.91,0.0,2313.8,0,0,91730
5207,0,1,1,0,24,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Credit card (automatic),40.65,933.3,1,74,32,0.0,3843,1,El Monte,1,0,DSL,34.079934,-118.046695,1,42.276,0,1,Offer C,30211,0,0,1,0,24,2,0.0,0.0,0.0,933.3,0,1,91731
5208,0,0,1,1,14,1,0,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),59.45,780.85,0,29,69,42.64,5723,0,El Monte,0,0,DSL,34.074492,-118.01462,1,59.45,2,4,Offer D,62660,1,0,1,0,14,0,0.0,596.96,0.0,780.85,1,1,91732
5209,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),109.95,7852.4,0,58,22,40.78,6258,0,South El Monte,0,1,Fiber Optic,34.04622,-118.053753,1,109.95,0,9,Offer A,45645,1,1,1,1,72,3,0.0,2936.16,0.0,7852.4,0,1,91733
5210,1,0,1,0,53,0,No phone service,DSL,0,1,1,1,One year,1,Electronic check,60.45,3184.25,1,61,14,0.0,5650,1,Rancho Cucamonga,1,1,DSL,34.245289,-117.642503,1,62.868,0,1,None,23079,1,1,1,1,53,2,446.0,0.0,0.0,3184.25,0,0,91737
5211,0,0,1,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.9,764.95,1,58,33,29.0,2656,1,Rancho Cucamonga,0,0,Fiber Optic,34.133809,-117.523724,1,88.296,0,1,None,12937,0,0,1,1,8,9,252.0,232.0,0.0,764.95,0,0,91739
5212,1,0,1,1,72,0,No phone service,DSL,1,1,0,0,Two year,0,Credit card (automatic),38.5,2763,0,25,82,0.0,4710,0,Glendora,1,1,DSL,34.119363,-117.85505900000001,1,38.5,3,8,Offer A,25135,0,0,1,0,72,0,2266.0,0.0,0.0,2763.0,1,0,91740
5213,0,1,1,0,17,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,92.55,1614.7,0,77,20,3.83,3689,0,Glendora,0,0,Fiber Optic,34.14649,-117.84981499999999,1,92.55,0,9,None,24973,0,0,1,0,17,0,32.29,65.11,0.0,1614.7,0,1,91741
5214,0,0,1,1,2,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),73.55,145.4,1,27,65,8.5,5799,1,La Puente,0,0,Cable,34.031441,-117.93643600000001,1,76.492,0,1,None,84965,0,1,1,1,2,1,9.45,17.0,0.0,145.4,1,1,91744
5215,0,0,1,0,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.15,156.25,1,24,0,11.35,4785,1,Hacienda Heights,0,0,NA,33.998471,-117.973758,1,20.15,0,1,None,53686,0,0,1,0,8,3,0.0,90.8,0.0,156.25,1,0,91745
5216,0,0,1,0,48,0,No phone service,DSL,0,1,0,0,One year,0,Mailed check,34.7,1604.5,1,31,24,0.0,5995,1,La Puente,1,0,Cable,34.038983,-117.991372,1,36.088,0,1,None,30802,0,3,1,0,48,1,385.0,0.0,0.0,1604.5,0,0,91746
5217,0,0,0,0,10,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,24.5,270.15,0,51,0,17.01,5594,0,Rowland Heights,0,0,NA,33.976753,-117.89736699999999,0,24.5,0,0,Offer D,46342,0,0,0,0,10,2,0.0,170.10000000000005,0.0,270.15,0,0,91748
5218,1,0,1,1,0,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.7, ,0,38,0,46.23,4890,0,La Verne,0,1,NA,34.144703,-117.770299,1,19.7,2,5,Offer E,35530,0,0,1,0,10,1,0.0,462.3,0.0,197.54,0,0,91750
5219,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.6,20.6,0,55,0,1.48,5370,0,Mira Loma,0,1,NA,33.999992,-117.535395,0,20.6,0,0,Offer E,18980,0,0,0,0,1,1,0.0,1.48,0.0,20.6,0,0,91752
5220,0,0,0,0,29,1,0,DSL,1,0,0,0,One year,0,Credit card (automatic),58.0,1734.5,0,42,25,14.46,2810,0,Monterey Park,1,0,Cable,34.050321999999994,-118.14703700000001,0,58.0,0,0,None,33280,1,0,0,0,29,2,434.0,419.34,0.0,1734.5,0,0,91754
5221,0,1,1,1,65,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,107.45,7047.5,0,65,26,19.58,6211,0,Monterey Park,1,0,Cable,34.049172,-118.115022,1,107.45,3,7,Offer B,26933,0,0,1,1,65,2,1832.0,1272.6999999999996,0.0,7047.5,0,0,91755
5222,0,0,0,0,8,1,1,DSL,1,1,0,0,Month-to-month,1,Bank transfer (automatic),65.5,573.15,0,37,28,8.73,3033,0,Mt Baldy,1,0,Fiber Optic,34.231318,-117.66203200000001,0,65.5,0,0,Offer E,47,0,0,0,0,8,1,160.0,69.84,0.0,573.15,0,0,91759
5223,1,0,1,0,61,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.45,1538.6,0,48,0,11.53,6015,0,Ontario,0,1,NA,34.035602000000004,-117.591528,1,25.45,0,2,Offer B,56280,0,1,1,0,61,1,0.0,703.3299999999998,0.0,1538.6,0,0,91761
5224,0,1,0,0,45,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),100.15,4459.8,0,68,20,6.9,2636,0,Ontario,1,0,Cable,34.057256,-117.667677,0,100.15,0,0,Offer B,54254,0,0,0,0,45,2,0.0,310.5,0.0,4459.8,0,1,91762
5225,1,0,1,1,72,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),104.45,7459,0,35,12,17.49,4750,0,Montclair,1,1,Fiber Optic,34.072121,-117.698319,1,104.45,1,5,Offer A,34447,0,0,1,1,72,1,89.51,1259.28,0.0,7459.0,0,1,91763
5226,1,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,21.15,306.05,0,50,0,33.9,5209,0,Ontario,0,1,NA,34.074087,-117.60561799999999,1,21.15,2,8,Offer D,49474,0,0,1,0,12,2,0.0,406.8,0.0,306.05,0,0,91764
5227,1,0,0,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,96.2,639.7,0,22,48,45.93,4329,0,Diamond Bar,0,1,Fiber Optic,33.992416,-117.807874,0,96.2,0,0,None,46532,0,0,0,1,7,0,307.0,321.51,0.0,639.7,1,0,91765
5228,1,0,0,0,9,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.4,348.15,0,19,26,38.65,5457,0,Pomona,0,1,Fiber Optic,34.042286,-117.756106,0,44.4,0,0,Offer E,69974,0,0,0,0,9,0,0.0,347.85,0.0,348.15,1,1,91766
5229,0,1,1,0,43,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,107.55,4533.9,1,80,20,13.84,4423,1,Pomona,1,0,Cable,34.083086,-117.737997,1,111.852,0,1,None,46626,1,4,1,0,43,4,907.0,595.12,0.0,4533.9,0,0,91767
5230,1,0,1,1,58,1,1,Fiber optic,0,0,0,1,Two year,0,Bank transfer (automatic),94.35,5563.65,0,54,23,5.01,4777,0,Pomona,1,1,DSL,34.067932,-117.785168,1,94.35,2,2,Offer B,36057,1,0,1,1,58,0,1280.0,290.58,0.0,5563.65,0,0,91768
5231,1,1,1,0,16,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.75,1587.55,1,69,8,15.16,3392,1,Rosemead,1,1,DSL,34.065108,-118.08279099999999,1,102.7,0,1,None,61623,0,2,1,0,16,2,127.0,242.56,0.0,1587.55,0,0,91770
5232,1,0,1,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.3,40.25,0,37,0,7.27,5113,0,San Dimas,0,1,NA,34.102119,-117.815532,1,20.3,2,5,Offer E,33878,0,0,1,0,2,0,0.0,14.54,0.0,40.25,0,0,91773
5233,0,0,1,0,8,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,101.15,842.9,1,47,7,16.88,2750,1,San Diego,1,0,DSL,32.787836,-117.232376,1,105.196,0,1,None,46086,0,0,1,1,8,0,59.0,135.04,0.0,842.9,0,0,92109
5234,0,0,1,0,40,1,1,Fiber optic,1,0,1,1,One year,0,Bank transfer (automatic),105.75,4228.55,0,24,76,22.2,4078,0,San Gabriel,1,0,Cable,34.089927,-118.09564499999999,1,105.75,0,5,Offer B,38041,0,0,1,1,40,0,0.0,888.0,0.0,4228.55,1,1,91776
5235,1,0,0,0,9,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,81.15,784.45,0,43,6,34.34,4544,0,Temple City,0,1,Fiber Optic,34.101608,-118.055848,0,81.15,0,0,Offer E,32718,0,0,0,0,9,0,0.0,309.06000000000006,0.0,784.45,0,1,91780
5236,1,0,0,0,41,1,0,Fiber optic,0,1,1,0,One year,1,Electronic check,89.55,3729.75,0,62,15,45.22,5549,0,Upland,0,1,Cable,34.141146,-117.65558300000001,0,89.55,0,0,Offer B,23331,1,0,0,0,41,3,0.0,1854.02,0.0,3729.75,0,1,91784
5237,0,0,0,0,26,1,0,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),54.75,1406.9,0,27,42,39.84,4020,0,Upland,1,0,Fiber Optic,34.105493,-117.66093400000001,0,54.75,0,0,None,48827,0,0,0,0,26,0,0.0,1035.84,0.0,1406.9,1,1,91786
5238,0,0,1,0,33,1,0,DSL,0,1,0,0,One year,1,Credit card (automatic),53.75,1857.3,0,27,59,15.45,3160,0,Walnut,0,0,Fiber Optic,34.018353999999995,-117.85491999999999,1,53.75,0,1,None,45118,1,0,1,0,33,0,1096.0,509.85,0.0,1857.3,1,0,91789
5239,1,0,1,1,68,1,0,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),105.75,7322.5,0,56,17,8.88,4437,0,West Covina,1,1,DSL,34.066964,-117.93700700000001,1,105.75,2,9,None,44099,1,0,1,1,68,1,0.0,603.84,0.0,7322.5,0,1,91790
5240,0,1,1,0,65,1,0,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),105.85,6725.5,0,65,9,36.49,4872,0,West Covina,1,0,DSL,34.061634000000005,-117.893169,1,105.85,0,10,Offer B,30458,1,0,1,1,65,0,60.53,2371.85,0.0,6725.5,0,1,91791
5241,1,0,0,0,55,1,0,DSL,0,1,0,1,One year,1,Electronic check,64.2,3627.3,0,47,26,27.65,5151,0,West Covina,0,1,DSL,34.024405,-117.89872199999999,0,64.2,0,0,Offer B,31622,1,0,0,1,55,3,943.0,1520.75,0.0,3627.3,0,0,91792
5242,1,0,0,0,20,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,88.7,1761.45,1,20,65,5.54,4115,1,San Diego,1,1,Cable,32.787836,-117.232376,0,92.24799999999999,0,0,Offer D,46086,0,0,0,0,20,2,1145.0,110.8,0.0,1761.45,1,0,92109
5243,1,0,0,0,19,1,0,Fiber optic,0,0,0,1,One year,1,Credit card (automatic),87.7,1725.95,0,49,2,43.11,4446,0,Alhambra,0,1,Fiber Optic,34.074736,-118.145959,0,87.7,0,0,Offer D,30635,1,0,0,1,19,0,35.0,819.09,0.0,1725.95,0,0,91803
5244,0,0,0,0,45,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),89.3,4192.15,0,42,8,13.82,5470,0,Alpine,1,0,Cable,32.827184,-116.70372900000001,0,89.3,0,0,Offer B,16486,0,0,0,1,45,0,0.0,621.9,0.0,4192.15,0,1,91901
5245,0,0,1,1,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.15,1411.2,0,32,0,26.85,5219,0,Bonita,0,0,NA,32.671170000000004,-117.00232,1,20.15,1,0,None,17389,0,0,0,0,70,0,0.0,1879.5,0.0,1411.2,0,0,91902
5246,0,0,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.75,164.5,1,44,18,8.32,5172,1,San Diego,0,0,Cable,32.787836,-117.232376,0,82.94,0,0,None,46086,0,0,0,0,2,2,30.0,16.64,0.0,164.5,0,0,92109
5247,0,0,0,0,27,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,94.55,2724.6,1,48,7,11.09,4464,1,San Diego,0,0,DSL,32.787836,-117.232376,0,98.33200000000001,0,0,None,46086,0,0,0,1,27,4,191.0,299.43,0.0,2724.6,0,0,92109
5248,0,0,1,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Electronic check,20.05,264.55,0,60,0,40.34,5453,0,Chula Vista,0,0,NA,32.636792,-117.05498899999999,1,20.05,0,10,Offer D,74025,0,0,1,0,12,0,0.0,484.08,0.0,264.55,0,0,91910
5249,1,0,0,1,72,0,No phone service,DSL,1,1,1,1,Two year,0,Credit card (automatic),67.2,4671.7,0,20,71,0.0,5592,0,Chula Vista,1,1,DSL,32.607964,-117.059459,0,67.2,3,0,None,71126,1,0,0,1,72,0,3317.0,0.0,0.0,4671.7,1,0,91911
5250,1,0,0,0,12,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,94.55,1173.55,0,38,8,13.88,5674,0,Chula Vista,0,1,DSL,32.64164,-116.985026,0,94.55,0,0,Offer D,12884,0,0,0,1,12,1,0.0,166.56,0.0,1173.55,0,1,91913
5251,0,1,0,0,5,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.05,318.5,1,71,12,30.05,3368,1,San Diego,0,0,Fiber Optic,32.787836,-117.232376,0,71.812,0,0,None,46086,0,1,0,0,5,2,38.0,150.25,0.0,318.5,0,0,92109
5252,1,1,1,0,71,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,107.5,7713.55,0,68,19,30.59,5775,0,Chula Vista,1,1,Cable,32.605012,-116.97595,1,107.5,0,7,None,9278,0,0,1,0,71,1,0.0,2171.89,0.0,7713.55,0,1,91915
5253,1,1,0,0,35,1,0,DSL,0,0,1,1,One year,1,Electronic check,73.0,2471.25,0,79,18,3.04,2715,0,Descanso,1,1,Fiber Optic,32.912664,-116.63538700000001,0,73.0,0,0,None,1587,1,0,0,0,35,2,44.48,106.4,0.0,2471.25,0,1,91916
5254,1,0,1,1,70,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),114.75,7842.3,0,54,75,39.06,5035,0,Dulzura,1,1,Fiber Optic,32.622999,-116.687855,1,114.75,3,10,None,727,1,0,1,1,70,0,5882.0,2734.2000000000007,0.0,7842.3,0,0,91917
5255,0,0,0,0,31,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.05,2227.8,0,30,59,38.78,2421,0,Guatay,0,0,Fiber Optic,32.857946000000005,-116.561917,0,76.05,0,0,None,796,0,1,0,0,31,2,131.44,1202.18,0.0,2227.8,0,1,91931
5256,1,0,1,1,52,1,1,Fiber optic,0,0,0,1,Two year,1,Bank transfer (automatic),96.25,4990.25,1,63,29,46.59,4751,1,San Diego,1,1,Cable,32.787836,-117.232376,1,100.1,0,1,None,46086,1,0,1,1,52,5,1447.0,2422.6800000000007,0.0,4990.25,0,0,92109
5257,1,1,0,0,37,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.1,3744.05,1,73,21,38.06,4424,1,San Diego,1,1,DSL,32.787836,-117.232376,0,105.144,0,0,Offer C,46086,0,0,0,0,37,2,0.0,1408.22,0.0,3744.05,0,1,92109
5258,1,0,0,0,69,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),104.7,7220.35,1,52,3,20.44,6350,1,San Diego,0,1,Fiber Optic,32.787836,-117.232376,0,108.88799999999999,0,0,Offer A,46086,1,0,0,1,69,3,0.0,1410.36,0.0,7220.35,0,1,92109
5259,1,1,1,0,30,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,77.9,2351.45,0,65,19,2.86,2009,0,La Mesa,0,1,DSL,32.759327,-116.99726000000001,1,77.9,0,1,None,44652,0,0,1,0,30,0,447.0,85.8,0.0,2351.45,0,0,91941
5260,0,0,0,0,33,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,90.65,2989.6,0,26,85,16.76,4460,0,La Mesa,0,0,DSL,32.782501,-117.01611000000001,0,90.65,0,0,None,24005,0,0,0,1,33,0,0.0,553.08,0.0,2989.6,1,1,91942
5261,1,1,1,0,54,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,110.45,6077.75,0,77,16,32.56,4425,0,Lemon Grove,1,1,DSL,32.733564,-117.03371299999999,1,110.45,0,5,Offer B,24961,1,0,1,0,54,0,972.0,1758.2400000000002,0.0,6077.75,0,0,91945
5262,0,0,0,0,59,1,1,DSL,1,0,0,1,One year,0,Bank transfer (automatic),68.7,4070.95,0,62,9,28.32,4244,0,Mount Laguna,0,0,Cable,32.830852,-116.444601,0,68.7,0,0,Offer B,81,1,0,0,1,59,1,0.0,1670.88,0.0,4070.95,0,1,91948
5263,1,1,0,0,55,0,No phone service,DSL,1,1,1,0,Month-to-month,1,Electronic check,44.85,2479.05,0,77,30,0.0,5829,0,National City,0,1,Cable,32.67102,-117.095235,0,44.85,0,0,Offer B,62355,0,0,0,0,55,0,0.0,0.0,0.0,2479.05,0,1,91950
5264,1,1,1,0,69,0,No phone service,DSL,0,0,0,0,One year,1,Credit card (automatic),29.8,2134.3,0,69,13,0.0,5681,0,Pine Valley,1,1,DSL,32.800671,-116.48336299999998,1,29.8,0,7,None,1604,0,0,1,0,69,0,0.0,0.0,0.0,2134.3,0,1,91962
5265,0,0,0,0,66,1,1,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),88.9,6000.1,0,33,15,31.93,5868,0,Potrero,0,0,Fiber Optic,32.619465000000005,-116.59360500000001,0,88.9,0,0,None,905,0,0,0,0,66,0,90.0,2107.38,0.0,6000.1,0,1,91963
5266,1,0,1,1,37,1,0,DSL,1,0,0,0,One year,1,Mailed check,58.75,2203.1,0,28,76,35.67,3483,0,Spring Valley,1,1,Cable,32.726627,-116.99460800000001,1,58.75,3,1,None,56100,1,0,1,0,37,3,0.0,1319.79,0.0,2203.1,1,1,91977
5267,1,1,1,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.85,183.15,0,79,0,22.79,5601,0,Spring Valley,0,1,NA,32.730264,-116.95096299999999,1,19.85,0,3,None,7863,0,0,1,0,9,1,0.0,205.11,0.0,183.15,0,0,91978
5268,1,0,1,1,69,1,1,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),86.9,6194.1,0,47,53,26.35,4667,0,Tecate,1,1,Cable,32.587557000000004,-116.636816,1,86.9,3,9,None,91,1,0,1,1,69,1,0.0,1818.15,0.0,6194.1,0,1,91980
5269,1,0,0,0,10,1,0,DSL,0,1,1,0,Month-to-month,1,Mailed check,59.65,638.95,0,36,25,1.48,2385,0,Bonsall,0,1,Fiber Optic,33.290907000000004,-117.202895,0,59.65,0,0,Offer D,3849,0,0,0,0,10,2,0.0,14.8,0.0,638.95,0,1,92003
5270,1,0,0,1,40,1,0,DSL,1,1,0,0,Month-to-month,1,Mailed check,55.25,2139.2,1,20,84,8.08,2810,1,San Diego,0,1,DSL,32.787836,-117.232376,0,57.46,1,0,None,46086,0,0,0,0,40,2,1797.0,323.2,0.0,2139.2,1,0,92109
5271,1,0,0,1,13,1,0,DSL,0,0,1,1,Month-to-month,0,Credit card (automatic),66.4,831.75,0,50,17,30.19,3660,0,Cardiff By The Sea,0,1,DSL,33.015865999999995,-117.272254,0,66.4,1,0,Offer D,10375,0,0,0,1,13,0,141.0,392.47,0.0,831.75,0,0,92007
5272,0,0,0,0,6,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,90.1,521.3,1,53,3,1.15,5656,1,San Diego,0,0,Fiber Optic,32.787836,-117.232376,0,93.704,0,0,None,46086,0,0,0,0,6,0,16.0,6.9,0.0,521.3,0,0,92109
5273,0,0,1,1,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.15,1337.5,0,64,0,11.47,4554,0,Carlsbad,0,0,NA,33.098017999999996,-117.25820300000001,1,20.15,3,6,None,43161,0,0,1,0,69,1,0.0,791.4300000000002,0.0,1337.5,0,0,92009
5274,0,1,1,0,66,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),108.1,7181.95,0,73,23,6.94,5360,0,Del Mar,1,0,Fiber Optic,32.948262,-117.25608600000001,1,108.1,0,3,None,13945,1,0,1,1,66,0,0.0,458.04,0.0,7181.95,0,1,92014
5275,1,0,0,0,11,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,53.75,608,1,60,14,15.03,3407,1,San Diego,1,1,Cable,32.787836,-117.232376,0,55.9,0,0,Offer D,46086,0,0,0,0,11,2,85.0,165.32999999999996,0.0,608.0,0,0,92109
5276,1,0,1,1,46,1,0,DSL,1,0,0,0,One year,0,Mailed check,56.9,2560.1,0,52,15,38.45,4258,0,El Cajon,1,1,Cable,32.79697,-116.969082,1,56.9,2,9,Offer B,55277,1,0,1,0,46,2,384.0,1768.7,0.0,2560.1,0,0,92020
5277,0,0,0,0,6,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,89.3,577.6,1,43,24,2.6,5800,1,San Diego,0,0,Cable,32.787836,-117.232376,0,92.87200000000001,0,0,None,46086,0,0,0,1,6,4,0.0,15.6,0.0,577.6,0,1,92109
5278,0,0,1,1,56,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Mailed check,109.6,5953,0,36,11,13.94,5012,0,Encinitas,1,0,Fiber Optic,33.054579,-117.25665,1,109.6,2,5,Offer B,47126,1,0,1,1,56,1,0.0,780.64,0.0,5953.0,0,1,92024
5279,1,0,1,1,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.15,1790.15,0,28,0,1.22,5114,0,Escondido,0,1,NA,33.081478000000004,-117.03381399999999,1,25.15,3,0,None,49281,0,0,0,0,70,0,0.0,85.39999999999998,0.0,1790.15,1,0,92025
5280,0,0,1,1,33,1,1,DSL,0,0,1,1,One year,1,Electronic check,79.15,2531.4,0,47,18,31.59,3555,0,Escondido,1,0,Fiber Optic,33.21846,-117.11691599999999,1,79.15,2,2,None,43436,1,0,1,1,33,0,45.57,1042.47,0.0,2531.4,0,1,92026
5281,0,0,1,1,72,1,1,DSL,1,1,0,0,Two year,0,Credit card (automatic),66.75,4760.3,0,56,27,22.62,6063,0,Escondido,0,0,Cable,33.141265000000004,-116.967221,1,66.75,3,8,None,48690,1,0,1,0,72,1,128.53,1628.64,0.0,4760.3,0,1,92027
5282,0,0,1,0,3,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.2,292.85,1,21,46,23.26,4176,1,San Diego,0,0,Fiber Optic,32.787836,-117.232376,1,99.008,0,5,None,46086,0,1,1,1,3,1,135.0,69.78,0.0,292.85,1,0,92109
5283,0,0,0,1,19,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,48.8,953.65,0,59,26,4.03,3749,0,Escondido,0,0,DSL,33.079834000000005,-117.134275,0,48.8,2,0,Offer D,17944,1,0,0,0,19,3,0.0,76.57000000000002,0.0,953.65,0,1,92029
5284,0,1,0,0,5,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Electronic check,45.7,198,1,79,16,0.0,3561,1,San Diego,0,0,Cable,32.787836,-117.232376,0,47.52800000000001,0,0,None,46086,0,2,0,0,5,3,32.0,0.0,0.0,198.0,0,0,92109
5285,0,0,1,0,71,1,0,DSL,0,1,1,1,Two year,1,Credit card (automatic),80.7,5705.05,0,48,27,43.61,5617,0,La Jolla,1,0,Fiber Optic,32.853743,-117.25034,1,80.7,0,8,None,42617,1,0,1,1,71,1,1540.0,3096.31,0.0,5705.05,0,0,92037
5286,1,0,1,0,8,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,74.5,609.9,1,51,25,47.91,3683,1,San Diego,0,1,Cable,32.787836,-117.232376,1,77.48,0,1,None,46086,0,0,1,0,8,2,152.0,383.28,0.0,609.9,0,0,92109
5287,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.55,20.55,0,29,0,7.32,4801,0,Oceanside,0,1,NA,33.351059,-117.420557,0,20.55,0,0,Offer E,98239,0,0,0,0,1,2,0.0,7.32,0.0,20.55,1,0,92054
5288,0,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.65,79.65,1,57,6,22.48,2119,1,San Diego,0,0,DSL,32.787836,-117.232376,0,82.83600000000001,0,0,None,46086,0,2,0,0,1,1,0.0,22.48,0.0,79.65,0,0,92109
5289,0,0,0,0,61,1,1,Fiber optic,1,1,1,1,One year,1,Mailed check,115.1,6993.65,0,58,7,5.55,4785,0,Oceanside,1,0,Cable,33.254497,-117.28587900000001,0,115.1,0,0,Offer B,46893,1,0,0,1,61,2,490.0,338.55,0.0,6993.65,0,0,92057
5290,0,0,1,1,71,0,No phone service,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),59.7,4122.65,0,44,19,0.0,6420,0,Pala,0,0,Cable,33.384345,-117.07261899999999,1,59.7,1,6,Offer A,1831,1,0,1,1,71,0,0.0,0.0,0.0,4122.65,0,1,92059
5291,0,0,1,0,68,1,1,Fiber optic,0,1,0,0,One year,0,Credit card (automatic),86.45,5762.95,0,48,15,9.76,4480,0,Palomar Mountain,1,0,Fiber Optic,33.309852,-116.82309099999999,1,86.45,0,5,Offer A,234,0,0,1,0,68,2,0.0,663.68,0.0,5762.95,0,1,92060
5292,1,0,0,0,46,0,No phone service,DSL,0,0,0,0,One year,0,Credit card (automatic),33.7,1537.85,0,35,18,0.0,3007,0,Pauma Valley,1,1,Fiber Optic,33.313828,-116.940501,0,33.7,0,0,Offer B,2615,1,1,0,0,46,1,277.0,0.0,0.0,1537.85,0,0,92061
5293,1,0,0,0,33,1,1,Fiber optic,1,0,0,0,One year,0,Bank transfer (automatic),80.1,2603.3,0,29,48,25.71,3957,0,Poway,0,1,Cable,32.984395,-117.01345400000001,0,80.1,0,0,None,47969,0,0,0,0,33,0,124.96,848.4300000000002,0.0,2603.3,1,1,92064
5294,0,0,1,1,53,1,1,Fiber optic,1,1,0,1,Two year,1,Bank transfer (automatic),104.05,5566.4,0,64,17,28.36,4190,0,Ramona,1,0,Fiber Optic,33.044540999999995,-116.833922,1,104.05,1,1,Offer B,33104,1,0,1,1,53,1,0.0,1503.08,0.0,5566.4,0,1,92065
5295,0,1,1,0,50,1,1,Fiber optic,1,1,1,1,Month-to-month,0,Bank transfer (automatic),108.75,5431.9,0,70,2,9.18,5211,0,Ranchita,1,0,Fiber Optic,33.215251,-116.53633,1,108.75,0,1,Offer B,339,0,0,1,1,50,0,109.0,459.0,0.0,5431.9,0,0,92066
5296,0,0,0,0,57,0,No phone service,DSL,1,0,0,0,One year,1,Credit card (automatic),41.1,2258.25,0,44,24,0.0,5281,0,Rancho Santa Fe,1,0,Fiber Optic,33.012751,-117.200617,0,41.1,0,0,None,7615,1,0,0,0,57,2,542.0,0.0,0.0,2258.25,0,0,92067
5297,0,0,1,1,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.35,1092.35,0,48,0,41.93,5646,0,San Marcos,0,0,NA,33.162624,-117.17086299999998,1,20.35,4,1,None,52664,0,0,1,0,54,1,0.0,2264.22,0.0,1092.35,0,0,92069
5298,0,1,1,0,60,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.9,6401.25,0,71,25,36.71,5084,0,Santa Ysabel,1,0,DSL,33.174725,-116.743329,1,105.9,0,1,Offer B,1143,0,0,1,1,60,1,1600.0,2202.6,0.0,6401.25,0,0,92070
5299,0,1,1,0,28,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),101.3,2812.2,1,67,22,16.43,4994,1,San Diego,0,0,Cable,32.787836,-117.232376,1,105.352,0,1,Offer C,46086,1,0,1,0,28,3,619.0,460.04,0.0,2812.2,0,0,92109
5300,0,0,1,1,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,80.05,80.05,1,53,8,39.79,2943,1,San Diego,0,0,Fiber Optic,32.787836,-117.232376,1,83.25200000000001,0,1,None,46086,0,1,1,0,1,2,0.0,39.79,0.0,80.05,0,0,92109
5301,1,0,1,1,29,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.2,2698.35,1,25,53,4.0,5292,1,San Diego,1,1,DSL,32.787836,-117.232376,1,92.76799999999999,0,1,None,46086,0,0,1,1,29,0,0.0,116.0,0.0,2698.35,1,1,92109
5302,0,0,1,1,10,1,0,DSL,0,1,0,1,Month-to-month,1,Electronic check,65.5,616.9,0,59,22,25.89,3137,0,Valley Center,0,0,Fiber Optic,33.252829999999996,-116.986079,1,65.5,1,1,Offer D,14575,1,0,1,1,10,2,136.0,258.9,0.0,616.9,0,0,92082
5303,1,0,0,1,43,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Electronic check,40.45,1912.85,0,41,25,0.0,3176,0,Vista,1,1,Fiber Optic,33.17494,-117.24276100000002,0,40.45,2,0,None,62036,0,0,0,0,43,0,0.0,0.0,0.0,1912.85,0,1,92083
5304,1,1,1,0,13,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),70.45,849.1,0,78,26,36.57,5225,0,Vista,0,1,Fiber Optic,33.22784,-117.200024,1,70.45,0,1,None,44692,0,1,1,0,13,2,22.08,475.41,0.0,849.1,0,1,92084
5305,0,0,1,0,43,1,0,DSL,1,0,1,1,Two year,1,Electronic check,78.8,3460.3,0,42,27,38.53,3972,0,Warner Springs,1,0,Fiber Optic,33.323705,-116.626907,1,78.8,0,1,None,1205,1,1,1,1,43,2,934.0,1656.79,24.9,3460.3,0,0,92086
5306,1,0,1,1,19,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,83.65,1465.75,1,59,28,14.09,3427,1,San Diego,0,1,Cable,32.787836,-117.232376,1,86.99600000000002,0,1,None,46086,0,0,1,1,19,0,410.0,267.71,0.0,1465.75,0,0,92109
5307,1,0,1,1,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,90.1,90.1,0,20,59,24.33,4142,0,San Diego,0,1,DSL,32.725229999999996,-117.171346,1,90.1,3,1,None,27505,0,0,1,1,1,0,0.0,24.33,0.0,90.1,1,1,92101
5308,0,0,0,0,69,1,0,DSL,1,0,1,1,Two year,1,Credit card (automatic),82.45,5555.3,0,46,22,25.73,4631,0,San Diego,1,0,DSL,32.716007,-117.11746200000002,0,82.45,0,0,Offer A,47140,1,0,0,1,69,1,122.22,1775.37,15.38,5555.3,0,1,92102
5309,0,0,1,0,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.25,1278.8,0,64,0,10.94,5974,0,San Diego,0,0,NA,32.747484,-117.166877,1,20.25,0,1,None,30202,0,1,1,0,61,1,0.0,667.3399999999998,5.15,1278.8,0,0,92103
5310,1,0,1,0,43,1,1,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),66.25,2907.35,0,42,17,26.1,2168,0,San Diego,0,1,Cable,32.741499,-117.12740900000001,1,66.25,0,1,None,47689,1,0,1,0,43,2,0.0,1122.3,6.41,2907.35,0,1,92104
5311,0,0,1,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.5,146.3,1,62,0,31.7,5579,1,San Diego,0,0,NA,32.787836,-117.232376,1,19.5,0,1,None,46086,0,0,1,0,6,3,0.0,190.2,0.0,146.3,0,0,92109
5312,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,51.25,51.25,1,58,4,6.44,2180,1,San Diego,0,1,Fiber Optic,32.787836,-117.232376,0,53.3,0,0,None,46086,1,0,0,0,1,0,0.0,6.44,0.0,51.25,0,0,92109
5313,1,0,1,0,56,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Mailed check,89.7,4952.95,0,43,14,3.79,5955,0,San Diego,0,1,Fiber Optic,32.741852,-117.243453,1,89.7,0,1,None,27959,0,0,1,1,56,0,693.0,212.24,41.66,4952.95,0,0,92107
5314,0,0,1,0,70,0,No phone service,DSL,1,1,1,1,Two year,0,Bank transfer (automatic),64.55,4504.9,0,21,46,0.0,4858,0,San Diego,1,0,Fiber Optic,32.774046000000006,-117.142454,1,64.55,0,5,Offer A,11650,1,0,1,1,70,0,2072.0,0.0,46.06,4504.9,1,0,92108
5315,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.6,45.6,1,31,26,11.73,3037,1,San Diego,0,1,Cable,32.787836,-117.232376,0,47.42400000000001,0,0,Offer E,46086,0,0,0,0,1,3,0.0,11.73,0.0,45.6,0,0,92109
5316,1,0,1,1,49,1,1,Fiber optic,0,1,1,0,One year,1,Electronic check,93.65,4520.15,0,27,59,36.08,5542,0,San Diego,1,1,DSL,32.76501,-117.19938,1,93.65,2,7,None,24169,0,0,1,0,49,1,2667.0,1767.9199999999996,33.13,4520.15,1,0,92110
5317,0,0,0,0,6,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),49.65,267.35,1,49,24,48.89,4248,1,San Diego,0,0,Cable,32.805518,-117.16905200000001,0,51.636,0,0,Offer E,46828,1,1,0,0,6,3,64.0,293.3400000000001,0.0,267.35,0,0,92111
5318,0,0,1,1,32,1,0,DSL,1,1,0,1,Two year,0,Mailed check,73.6,2316.85,0,26,59,19.76,4343,0,San Diego,1,0,DSL,32.697098,-117.11658700000001,1,73.6,1,1,None,47431,1,0,1,1,32,1,0.0,632.32,12.66,2316.85,1,1,92113
5319,0,1,1,0,72,1,1,Fiber optic,1,0,1,1,Two year,1,Mailed check,109.75,8075.35,0,73,22,35.04,6010,0,San Diego,1,0,Cable,32.707892,-117.05512,1,109.75,0,1,Offer A,66838,1,0,1,0,72,1,1777.0,2522.88,0.0,8075.35,0,0,92114
5320,1,0,0,1,37,1,0,DSL,1,1,0,0,Two year,0,Credit card (automatic),61.45,2302.35,0,45,27,49.99,5447,0,San Diego,0,1,Fiber Optic,32.762506,-117.07245,0,61.45,1,0,None,56887,1,0,0,0,37,0,622.0,1849.63,48.79,2302.35,0,0,92115
5321,0,0,1,0,69,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),106.4,7251.9,0,59,5,24.17,4328,0,San Diego,0,0,Cable,32.765299,-117.122565,1,106.4,0,9,Offer A,33083,1,0,1,1,69,0,36.26,1667.73,3.59,7251.9,0,1,92116
5322,0,0,1,0,26,1,0,DSL,0,1,1,1,Month-to-month,0,Bank transfer (automatic),81.9,2078.55,0,26,48,11.23,3350,0,San Diego,1,0,Fiber Optic,32.825086,-117.199424,1,81.9,0,7,None,51213,1,0,1,1,26,3,0.0,291.98,44.86,2078.55,1,1,92117
5323,0,0,1,1,58,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),105.2,6225.4,0,61,30,43.01,4605,0,Coronado,1,0,Fiber Optic,32.68674,-117.18661200000001,1,105.2,3,2,None,24093,0,0,1,1,58,2,0.0,2494.58,34.83,6225.4,0,1,92118
5324,1,0,0,0,24,1,1,DSL,0,0,0,0,One year,0,Bank transfer (automatic),54.6,1242.25,0,28,85,7.52,3398,0,San Diego,0,1,Fiber Optic,32.802959,-117.02709499999999,0,54.6,0,0,None,21866,1,0,0,0,24,1,105.59,180.48,28.42,1242.25,1,1,92119
5325,1,0,1,1,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,20.55,99.45,0,27,0,41.21,3629,0,San Diego,0,1,NA,32.807867,-117.060993,1,20.55,2,1,None,25569,0,0,1,0,5,1,0.0,206.05,0.0,99.45,1,0,92120
5326,1,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.0,288.05,1,59,0,31.14,4672,1,San Diego,0,1,NA,32.898613,-117.202937,1,20.0,3,1,None,4258,0,1,1,0,15,2,0.0,467.1,0.0,288.05,0,0,92121
5327,0,0,1,1,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.7,599.25,0,24,0,12.85,5045,0,San Diego,0,0,NA,32.85723,-117.209774,1,19.7,1,1,None,34902,0,0,1,0,30,0,0.0,385.5,49.79,599.25,1,0,92122
5328,0,0,1,0,55,1,1,DSL,1,1,0,0,One year,1,Credit card (automatic),66.05,3462.1,0,41,13,35.38,5501,0,San Diego,0,0,Fiber Optic,32.808814,-117.134694,1,66.05,0,0,None,25232,1,0,0,0,55,0,0.0,1945.9,44.53,3462.1,0,1,92123
5329,0,0,1,0,25,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Bank transfer (automatic),34.0,853,1,19,90,0.0,5024,1,San Diego,0,0,Cable,32.827238,-117.08928700000001,1,35.36,0,1,Offer C,30206,0,4,1,0,25,1,768.0,0.0,0.0,853.0,1,0,92124
5330,1,1,1,0,10,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Mailed check,92.5,934.1,1,72,33,11.12,2415,1,San Diego,1,1,DSL,32.886925,-117.152162,1,96.2,0,1,None,74232,1,0,1,0,10,2,0.0,111.2,0.0,934.1,0,1,92126
5331,1,0,1,1,44,0,No phone service,DSL,1,1,0,1,Two year,1,Credit card (automatic),54.05,2375.2,0,19,59,0.0,4896,0,San Diego,1,1,Fiber Optic,33.017518,-117.11845600000001,1,54.05,2,1,None,20046,1,0,1,1,44,1,0.0,0.0,47.45,2375.2,1,1,92127
5332,0,0,0,0,47,1,0,DSL,1,1,0,0,One year,1,Mailed check,58.9,2813.05,0,55,5,26.35,5774,0,San Diego,0,0,Fiber Optic,33.000269,-117.072093,0,58.9,0,0,None,42733,1,0,0,0,47,1,14.07,1238.45,0.0,2813.05,0,1,92128
5333,0,0,1,1,13,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,88.35,1222.8,1,52,11,17.83,3740,1,San Diego,0,0,DSL,32.886925,-117.152162,1,91.884,0,1,None,74232,0,0,1,1,13,4,135.0,231.79,0.0,1222.8,0,0,92126
5334,0,0,1,1,49,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),107.95,5293.2,1,38,11,6.45,5785,1,San Diego,1,0,DSL,32.886925,-117.152162,1,112.26799999999999,0,1,None,74232,1,0,1,1,49,6,0.0,316.05,0.0,5293.2,0,1,92126
5335,0,0,1,0,64,1,0,Fiber optic,1,0,1,1,One year,1,Mailed check,96.9,6314.35,0,31,21,19.22,5369,0,San Diego,0,0,DSL,32.89325,-117.08709099999999,1,96.9,0,10,None,29283,1,0,1,1,64,2,1326.0,1230.08,13.37,6314.35,0,0,92131
5336,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.1,19.1,0,61,0,44.22,2091,0,San Diego,0,1,NA,32.677716,-117.04766599999999,0,19.1,0,0,None,36351,0,0,0,0,1,3,0.0,44.22,0.0,19.1,0,0,92139
5337,1,0,0,0,20,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,50.0,1003.05,0,38,4,49.81,5741,0,San Diego,0,1,Cable,32.578103000000006,-117.012975,0,50.0,0,0,Offer D,68776,1,0,0,0,20,0,4.01,996.2,2.81,1003.05,0,1,92154
5338,0,0,1,0,37,0,No phone service,DSL,1,0,1,0,Two year,0,Electronic check,45.4,1593.1,0,23,27,0.0,4051,0,San Ysidro,0,0,Fiber Optic,32.555828000000005,-117.04007299999999,1,45.4,0,1,None,28488,1,1,1,0,37,2,0.0,0.0,44.13,1593.1,1,1,92173
5339,1,0,1,1,30,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,85.45,2509.95,0,63,19,21.72,3409,0,Indio,0,1,Fiber Optic,33.713891,-116.237257,1,85.45,2,9,None,56307,0,0,1,0,30,0,477.0,651.5999999999998,23.13,2509.95,0,0,92201
5340,0,0,0,0,38,1,1,DSL,1,1,1,1,One year,0,Bank transfer (automatic),84.1,3187.65,0,57,13,25.11,2604,0,Indio,1,0,DSL,33.752938,-116.23005500000001,0,84.1,0,0,None,2743,0,0,0,1,38,0,0.0,954.18,0.0,3187.65,0,1,92203
5341,0,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.45,74.45,1,75,18,39.61,4291,1,San Diego,0,0,DSL,32.886925,-117.152162,0,77.42800000000003,0,0,None,74232,0,0,0,0,1,0,0.0,39.61,0.0,74.45,0,0,92126
5342,0,0,0,0,37,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,64.75,2345.2,1,26,78,3.27,5554,1,San Diego,0,0,DSL,32.886925,-117.152162,0,67.34,0,0,Offer C,74232,0,2,0,1,37,2,1829.0,120.99,0.0,2345.2,1,0,92126
5343,0,0,1,0,52,0,No phone service,DSL,1,1,1,1,Two year,0,Credit card (automatic),66.25,3330.1,0,22,52,0.0,4275,0,Banning,1,0,Cable,33.936298,-116.849577,1,66.25,0,3,None,25859,1,0,1,1,52,0,1732.0,0.0,0.0,3330.1,1,0,92220
5344,1,0,0,1,71,1,0,DSL,1,1,1,0,Two year,1,Credit card (automatic),76.9,5522.7,0,20,52,4.76,4633,0,Beaumont,1,1,Fiber Optic,33.946982,-116.977672,0,76.9,3,0,Offer A,17721,1,0,0,0,71,0,0.0,337.96,0.0,5522.7,1,1,92223
5345,1,0,0,0,26,1,0,Fiber optic,0,1,1,0,Month-to-month,0,Electronic check,89.8,2335.3,1,49,28,6.24,3452,1,San Diego,1,1,Cable,32.886925,-117.152162,0,93.39200000000001,0,0,Offer C,74232,0,1,0,0,26,3,654.0,162.24,0.0,2335.3,0,0,92126
5346,1,0,0,0,66,1,1,DSL,1,1,0,1,Two year,1,Credit card (automatic),74.6,4798.4,0,56,11,45.57,4838,0,Brawley,1,1,Cable,33.03933,-115.19185700000001,0,74.6,0,0,Offer A,23394,0,0,0,1,66,1,0.0,3007.62,0.0,4798.4,0,1,92227
5347,1,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),116.95,8594.4,0,45,3,17.87,5949,0,Cabazon,1,1,Fiber Optic,33.929812,-116.76058,1,116.95,0,9,Offer A,2355,1,0,1,1,72,2,258.0,1286.64,0.0,8594.4,0,0,92230
5348,1,0,0,1,25,0,No phone service,DSL,1,0,1,0,One year,1,Credit card (automatic),40.65,970.55,0,56,18,0.0,5079,0,Calexico,0,1,DSL,32.690653999999995,-115.431225,0,40.65,2,0,None,27804,0,0,0,0,25,0,175.0,0.0,0.0,970.55,0,0,92231
5349,1,0,1,1,69,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.35,7665.8,0,24,27,37.97,6082,0,Calipatria,1,1,Fiber Optic,33.143826000000004,-115.49748500000001,1,114.35,3,7,Offer A,7857,1,0,1,1,69,1,0.0,2619.93,0.0,7665.8,1,1,92233
5350,1,0,1,1,53,1,1,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),69.7,3686.05,0,54,57,27.93,4975,0,Cathedral City,0,1,DSL,33.829583,-116.474131,1,69.7,3,9,None,43141,0,0,1,1,53,1,0.0,1480.29,0.0,3686.05,0,1,92234
5351,0,0,0,0,12,1,0,Fiber optic,0,0,1,1,One year,0,Mailed check,95.5,1115.15,1,61,18,34.81,3538,1,San Diego,1,0,Fiber Optic,32.886925,-117.152162,0,99.32,0,0,None,74232,0,2,0,1,12,8,0.0,417.72,0.0,1115.15,0,1,92126
5352,1,0,0,0,26,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.65,2537,0,26,76,37.0,4191,0,Desert Center,1,1,Fiber Optic,33.889604999999996,-115.25700900000001,0,98.65,0,0,None,964,1,0,0,1,26,2,0.0,962.0,0.0,2537.0,1,1,92239
5353,1,0,0,0,21,1,0,DSL,0,0,0,1,Month-to-month,0,Mailed check,61.65,1393.6,0,25,52,39.85,2926,0,Desert Hot Springs,1,1,Cable,33.948558,-116.516976,0,61.65,0,0,Offer D,22796,0,0,0,1,21,0,72.47,836.85,0.0,1393.6,1,1,92240
5354,0,0,0,1,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.35,89.35,0,38,19,5.36,2432,0,Desert Hot Springs,0,0,DSL,33.832799,-116.250973,0,89.35,1,0,None,5529,0,0,0,1,1,0,0.0,5.36,0.0,89.35,0,0,92241
5355,1,0,0,0,48,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,95.4,4445.3,0,28,46,4.15,4334,0,Earp,0,1,Cable,34.137741999999996,-114.36514,0,95.4,0,0,None,1564,1,1,0,1,48,2,2045.0,199.2,0.0,4445.3,1,0,92242
5356,0,0,1,0,26,0,No phone service,DSL,1,0,0,0,One year,0,Credit card (automatic),35.4,978.6,0,24,51,0.0,2519,0,El Centro,1,0,DSL,32.770393,-115.60915,1,35.4,0,4,None,43712,0,1,1,0,26,2,49.91,0.0,0.0,978.6,1,1,92243
5357,1,0,1,0,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.95,1258.15,0,39,0,30.14,5971,0,Heber,0,1,NA,32.730583,-115.50108300000001,1,19.95,0,7,None,3535,0,0,1,0,60,0,0.0,1808.4,0.0,1258.15,0,0,92249
5358,1,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.25,331.35,0,50,0,31.33,4769,0,Holtville,0,1,NA,32.811001,-115.15286499999999,0,19.25,0,0,Offer D,8062,0,0,0,0,18,0,0.0,563.9399999999998,0.0,331.35,0,0,92250
5359,0,1,0,0,10,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,29.65,291.4,1,76,22,0.0,5702,1,San Diego,0,0,Fiber Optic,32.886925,-117.152162,0,30.836,0,0,None,74232,1,1,0,0,10,4,64.0,0.0,0.0,291.4,0,0,92126
5360,1,0,1,1,5,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,84.5,453.75,1,64,9,36.88,5141,1,San Diego,1,1,Cable,32.886925,-117.152162,1,87.88000000000002,0,3,Offer E,74232,0,0,1,0,5,7,0.0,184.4,0.0,453.75,0,1,92126
5361,0,0,0,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.4,84.75,0,52,0,32.15,5602,0,La Quinta,0,0,NA,33.695532,-116.310571,0,20.4,1,0,None,23971,0,1,0,0,4,1,0.0,128.6,0.0,84.75,0,0,92253
5362,1,0,1,1,65,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.75,1715.1,0,52,0,36.5,6263,0,Mecca,0,1,NA,33.543834999999994,-115.99390600000001,1,24.75,2,4,None,8768,0,0,1,0,65,0,0.0,2372.5,0.0,1715.1,0,0,92254
5363,1,0,1,1,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.35,1715.15,0,63,0,10.46,6059,0,Morongo Valley,0,1,NA,34.097863000000004,-116.59456100000001,1,25.35,1,6,Offer A,3499,0,1,1,0,70,3,0.0,732.2,0.0,1715.15,0,0,92256
5364,1,0,0,0,18,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),90.7,1597.25,1,26,29,28.59,2931,1,San Diego,1,1,DSL,32.886925,-117.152162,0,94.32799999999999,0,0,None,74232,0,0,0,1,18,1,463.0,514.62,0.0,1597.25,1,0,92126
5365,1,0,0,1,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.0,1250.1,0,44,0,24.48,4402,0,North Palm Springs,0,1,NA,33.906496000000004,-116.569499,0,20.0,2,0,None,732,0,0,0,0,62,0,0.0,1517.76,0.0,1250.1,0,0,92258
5366,0,0,1,1,66,1,0,DSL,1,0,1,0,Two year,1,Electronic check,59.75,3996.8,0,58,16,8.39,5979,0,Ocotillo,0,0,Fiber Optic,32.698964000000004,-115.886656,1,59.75,2,9,Offer A,471,0,0,1,0,66,2,0.0,553.74,0.0,3996.8,0,1,92259
5367,0,0,1,1,65,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),82.5,5215.1,0,23,69,4.75,5314,0,Palm Desert,0,0,Fiber Optic,33.694501,-116.41271100000002,1,82.5,2,0,Offer B,29340,1,0,0,1,65,2,3598.0,308.75,0.0,5215.1,1,0,92260
5368,0,1,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,235.5,1,69,18,5.54,5165,1,San Diego,0,0,Fiber Optic,32.886925,-117.152162,0,73.112,0,0,None,74232,0,0,0,0,3,3,42.0,16.62,0.0,235.5,0,0,92126
5369,0,0,0,0,34,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,673.2,0,19,0,36.75,2864,0,Palm Springs,0,0,NA,33.745746000000004,-116.514215,0,20.35,0,0,None,18884,0,0,0,0,34,1,0.0,1249.5,0.0,673.2,1,0,92264
5370,1,0,1,1,16,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),90.8,1442.2,0,49,12,48.71,5560,0,Palo Verde,1,1,DSL,33.3249,-114.758334,1,90.8,2,8,Offer D,291,0,1,1,0,16,1,0.0,779.36,0.0,1442.2,0,1,92266
5371,0,0,0,0,54,1,1,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),103.95,5639.05,1,20,90,43.47,6117,1,San Diego,1,0,Cable,32.886925,-117.152162,0,108.10799999999999,0,0,None,74232,0,0,0,1,54,2,5075.0,2347.38,0.0,5639.05,1,0,92126
5372,0,1,0,0,50,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,104.95,5222.35,0,75,29,17.65,5570,0,Pioneertown,1,0,Fiber Optic,34.201108000000005,-116.593456,0,104.95,0,0,Offer B,354,1,0,0,0,50,0,0.0,882.4999999999999,0.0,5222.35,0,1,92268
5373,1,0,1,0,71,1,0,Fiber optic,0,1,1,1,Two year,1,Electronic check,105.25,7291.75,0,54,8,37.69,6319,0,Rancho Mirage,1,1,Cable,33.763678000000006,-116.429928,1,105.25,0,10,Offer A,12465,1,0,1,1,71,0,58.33,2675.99,0.0,7291.75,0,1,92270
5374,0,0,0,0,10,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.75,799.65,1,39,29,5.63,5578,1,San Diego,0,0,DSL,32.886925,-117.152162,0,77.74000000000002,0,0,None,74232,0,2,0,0,10,2,232.0,56.3,0.0,799.65,0,0,92126
5375,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.8,50.8,1,20,30,22.82,4535,1,San Diego,0,0,Fiber Optic,32.886925,-117.152162,0,52.832,0,0,None,74232,1,0,0,0,1,3,0.0,22.82,0.0,50.8,1,0,92126
5376,1,0,0,0,18,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,23.75,424.5,0,45,0,12.97,3076,0,Salton City,0,1,NA,33.28156,-115.955541,0,23.75,0,0,Offer D,799,0,0,0,0,18,0,0.0,233.46,0.0,424.5,0,0,92275
5377,1,0,0,0,4,1,0,DSL,0,0,1,0,Month-to-month,1,Electronic check,61.3,249.4,0,54,2,37.7,5281,0,Thousand Palms,0,1,Fiber Optic,33.849263,-116.382778,0,61.3,0,0,None,6242,1,0,0,0,4,0,0.0,150.8,0.0,249.4,0,1,92276
5378,0,0,1,1,58,1,1,DSL,1,0,1,0,Two year,0,Mailed check,75.8,4415.75,0,28,69,2.87,4292,0,Escondido,1,0,Fiber Optic,33.141265000000004,-116.967221,1,75.8,2,1,Offer B,48690,1,0,1,0,58,1,3047.0,166.46,0.0,4415.75,1,0,92027
5379,0,0,1,0,56,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,98.0,5270.6,0,33,11,37.5,4615,0,Twentynine Palms,0,0,Cable,34.457829,-116.13958899999999,1,98.0,0,10,Offer B,14104,0,0,1,1,56,1,580.0,2100.0,0.0,5270.6,0,0,92278
5380,1,0,0,0,2,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.25,144.55,1,42,33,39.03,5055,1,San Diego,0,1,DSL,32.886925,-117.152162,0,83.46000000000002,0,0,Offer E,74232,0,0,0,0,2,4,48.0,78.06,0.0,144.55,0,0,92126
5381,1,0,1,0,32,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,78.9,2447.95,1,62,12,22.57,5949,1,San Diego,1,1,Fiber Optic,32.886925,-117.152162,1,82.05600000000003,0,1,Offer C,74232,0,1,1,0,32,5,294.0,722.24,0.0,2447.95,0,0,92126
5382,1,0,1,1,56,0,No phone service,DSL,1,1,1,0,One year,1,Mailed check,52.0,2884.9,0,24,41,0.0,5845,0,White Water,0,1,DSL,33.972293,-116.654195,1,52.0,2,8,Offer B,805,1,0,1,0,56,1,1183.0,0.0,0.0,2884.9,1,0,92282
5383,1,0,0,0,36,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.75,3050.15,1,22,46,43.97,5272,1,San Diego,0,1,Cable,32.886925,-117.152162,0,88.14,0,0,Offer C,74232,0,1,0,1,36,4,0.0,1582.92,0.0,3050.15,1,1,92126
5384,0,0,0,0,4,1,1,DSL,0,0,1,0,Month-to-month,1,Mailed check,64.4,253,0,58,19,1.1,3334,0,Yucca Valley,0,0,Fiber Optic,34.159534,-116.42598400000001,0,64.4,0,0,None,20486,1,0,0,0,4,0,0.0,4.4,0.0,253.0,0,1,92284
5385,1,0,0,0,53,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Bank transfer (automatic),85.45,4517.25,1,38,32,16.43,4753,1,San Diego,0,1,Fiber Optic,32.886925,-117.152162,0,88.86800000000002,0,0,None,74232,0,0,0,0,53,0,0.0,870.79,0.0,4517.25,0,1,92126
5386,1,0,0,0,10,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),45.8,436.2,0,34,22,15.45,5586,0,Adelanto,0,1,Fiber Optic,34.667815000000004,-117.53618300000001,0,45.8,0,0,None,18980,0,2,0,0,10,1,9.6,154.5,0.0,436.2,0,1,92301
5387,1,0,0,0,4,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,30.5,118.4,0,52,22,0.0,3030,0,Amboy,0,1,Fiber Optic,34.559882,-115.63716399999998,0,30.5,0,0,None,42,1,0,0,0,4,1,2.6,0.0,0.0,118.4,0,1,92304
5388,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,19.9,1,46,0,45.77,5441,1,San Diego,0,1,NA,32.886925,-117.152162,1,19.9,1,4,Offer E,74232,0,0,1,0,1,1,0.0,45.77,0.0,19.9,0,0,92126
5389,0,0,1,0,51,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,69.15,3649.6,0,63,13,45.76,5187,0,Fallbrook,0,0,Fiber Optic,33.362575,-117.299644,1,69.15,0,1,Offer B,42239,0,0,1,0,51,1,474.0,2333.76,0.0,3649.6,0,0,92028
5390,1,1,0,0,12,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,99.45,1200.15,1,76,29,21.89,2819,1,San Diego,1,1,DSL,32.886925,-117.152162,0,103.428,0,0,None,74232,0,0,0,0,12,2,0.0,262.68,0.0,1200.15,0,1,92126
5391,0,0,0,0,6,0,No phone service,DSL,0,0,1,1,One year,1,Mailed check,49.25,255.6,0,29,48,0.0,2979,0,Baker,0,0,Fiber Optic,35.28952,-116.09221399999998,0,49.25,0,0,None,904,1,1,0,1,6,1,0.0,0.0,0.0,255.6,1,1,92309
5392,1,0,1,1,63,0,No phone service,DSL,0,1,0,0,Two year,0,Bank transfer (automatic),39.35,2395.05,0,45,16,0.0,5374,0,Fort Irwin,1,1,Cable,35.349241,-116.77028100000001,1,39.35,2,7,Offer B,9465,1,0,1,0,63,2,383.0,0.0,0.0,2395.05,0,0,92310
5393,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.6,70.6,1,48,25,27.12,4063,1,San Diego,0,0,Fiber Optic,32.886925,-117.152162,0,73.42399999999998,0,0,None,74232,0,0,0,0,1,3,0.0,27.12,0.0,70.6,0,0,92126
5394,0,0,1,0,48,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),105.1,5083.55,0,22,51,39.25,3109,0,Grand Terrace,0,0,Fiber Optic,34.029175,-117.30721100000001,1,105.1,0,4,Offer B,11024,1,0,1,1,48,1,0.0,1884.0,0.0,5083.55,1,1,92313
5395,0,0,0,0,5,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),81.0,389.6,1,61,25,20.2,3718,1,San Diego,0,0,DSL,32.886925,-117.152162,0,84.24000000000002,0,0,Offer E,74232,0,0,0,0,5,1,0.0,101.0,0.0,389.6,0,1,92126
5396,0,0,0,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Credit card (automatic),20.1,644.5,0,44,0,25.52,3726,0,Big Bear Lake,0,0,NA,34.242058,-116.89801999999999,0,20.1,1,0,None,5447,0,0,0,0,35,0,0.0,893.1999999999998,0.0,644.5,0,0,92315
5397,1,0,0,0,6,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,84.85,523.5,1,61,13,39.32,3420,1,San Diego,0,1,DSL,32.886925,-117.152162,0,88.244,0,0,Offer E,74232,0,3,0,0,6,4,68.0,235.92,0.0,523.5,0,0,92126
5398,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.75,39.3,0,58,0,1.97,4064,0,Calimesa,0,1,NA,33.982787,-117.057627,0,19.75,0,0,None,7334,0,0,0,0,2,0,0.0,3.94,0.0,39.3,0,0,92320
5399,0,0,0,0,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.75,989.05,0,63,0,37.95,4934,0,Cedar Glen,0,0,NA,34.255203,-117.17565400000001,0,19.75,0,0,Offer B,455,0,0,0,0,50,2,0.0,1897.5,0.0,989.05,0,0,92321
5400,0,0,0,0,33,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),70.4,2406.1,0,43,19,49.45,4860,0,Colton,0,0,Fiber Optic,34.030915,-117.273201,0,70.4,0,0,None,52202,0,0,0,0,33,0,0.0,1631.85,0.0,2406.1,0,1,92324
5401,1,0,0,0,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.45,638.55,0,59,0,34.57,2598,0,Crestline,0,1,NA,34.248061,-117.29028000000001,0,20.45,0,0,None,10484,0,0,0,0,31,1,0.0,1071.67,0.0,638.55,0,0,92325
5402,0,0,1,1,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.35,191.1,0,22,0,30.83,5352,0,Daggett,0,0,NA,34.875144,-116.821698,1,20.35,1,9,None,678,0,0,1,0,9,0,0.0,277.47,0.0,191.1,1,0,92327
5403,0,0,1,1,54,1,1,DSL,0,1,1,1,Month-to-month,1,Electronic check,86.2,4524.05,0,40,12,4.33,6275,0,Death Valley,1,0,Fiber Optic,36.27688,-117.033326,1,86.2,2,7,Offer B,443,1,0,1,1,54,3,0.0,233.82,0.0,4524.05,0,1,92328
5404,0,0,0,0,46,1,0,Fiber optic,1,1,1,0,One year,1,Credit card (automatic),95.65,4664.2,0,27,59,30.6,4727,0,Essex,1,0,DSL,34.9436,-115.287901,0,95.65,0,0,Offer B,115,0,0,0,0,46,0,2752.0,1407.6,0.0,4664.2,1,0,92332
5405,1,0,0,1,34,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,103.8,3470.8,0,35,16,4.28,5382,0,Fawnskin,0,1,Fiber Optic,34.274846000000004,-116.93758100000001,0,103.8,1,0,Offer C,414,0,0,0,1,34,1,555.0,145.52,0.0,3470.8,0,0,92333
5406,1,0,1,1,71,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,97.2,6910.3,0,28,69,39.09,4603,0,Fontana,0,1,Fiber Optic,34.087558,-117.464096,1,97.2,2,7,Offer A,82630,0,0,1,1,71,0,0.0,2775.390000000001,0.0,6910.3,1,1,92335
5407,0,0,1,1,63,1,0,DSL,1,1,0,0,Two year,0,Mailed check,63.55,4014.2,0,62,27,1.18,5733,0,Fontana,1,0,Fiber Optic,34.136367,-117.460803,1,63.55,2,6,Offer B,54586,1,0,1,0,63,2,1084.0,74.33999999999997,0.0,4014.2,0,0,92336
5408,0,0,0,0,51,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.95,1288,0,56,0,44.35,5458,0,Fontana,0,0,NA,34.049671000000004,-117.468896,0,24.95,0,0,Offer B,29847,0,1,0,0,51,3,0.0,2261.85,0.0,1288.0,0,0,92337
5409,0,1,0,0,26,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.15,2277.65,1,68,13,9.09,4074,1,San Diego,0,0,Cable,32.886925,-117.152162,0,92.716,0,0,Offer C,74232,0,0,0,0,26,4,0.0,236.34,0.0,2277.65,0,1,92126
5410,0,0,1,0,64,1,0,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),99.0,6375.8,0,35,11,35.92,5483,0,Forest Falls,1,0,Fiber Optic,34.067699,-116.90389099999999,1,99.0,0,7,Offer B,958,0,0,1,1,64,2,701.0,2298.88,0.0,6375.8,0,0,92339
5411,0,1,1,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.8,24.8,1,77,21,0.0,5377,1,San Diego,0,0,DSL,32.886925,-117.152162,1,25.791999999999998,0,1,None,74232,0,0,1,0,1,3,0.0,0.0,0.0,24.8,0,1,92126
5412,1,1,1,0,61,1,1,Fiber optic,0,1,0,0,One year,1,Bank transfer (automatic),85.55,5251.75,0,78,23,46.65,4845,0,Helendale,0,1,Fiber Optic,34.757783,-117.33997,1,85.55,0,5,Offer B,4948,1,0,1,0,61,0,0.0,2845.65,0.0,5251.75,0,1,92342
5413,0,0,0,0,15,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),94.0,1505.45,0,54,16,15.28,4521,0,Hesperia,1,0,Fiber Optic,34.361387,-117.33750900000001,0,94.0,0,0,None,68515,0,0,0,1,15,0,241.0,229.2,0.0,1505.45,0,0,92345
5414,1,0,0,0,64,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),105.65,6903.1,1,30,80,24.23,4870,1,San Diego,0,1,Fiber Optic,32.886925,-117.152162,0,109.876,0,0,None,74232,1,1,0,1,64,5,5522.0,1550.72,0.0,6903.1,0,0,92126
5415,0,0,0,0,18,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.3,913.3,0,40,20,38.32,5877,0,Hinkley,0,0,Fiber Optic,34.983808,-117.239306,0,50.3,0,0,None,1933,0,0,0,0,18,0,0.0,689.76,0.0,913.3,0,1,92347
5416,0,0,1,1,57,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,95.0,5535.8,0,35,22,42.18,6245,0,Lake Arrowhead,0,0,Fiber Optic,34.2565,-117.19335,1,95.0,2,3,Offer B,9793,0,0,1,1,57,0,0.0,2404.26,0.0,5535.8,0,1,92352
5417,1,0,1,1,14,1,0,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),61.4,815.55,0,20,59,10.74,3186,0,Loma Linda,0,1,DSL,34.049315,-117.255974,1,61.4,1,3,None,18068,0,0,1,1,14,0,481.0,150.36,0.0,815.55,1,0,92354
5418,1,1,0,0,18,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),80.55,1411.65,0,67,14,38.79,5137,0,Lucerne Valley,0,1,DSL,34.508417,-116.856103,0,80.55,0,0,None,5256,0,0,0,0,18,2,0.0,698.22,0.0,1411.65,0,1,92356
5419,0,1,1,0,72,1,1,Fiber optic,1,0,0,0,Two year,0,Bank transfer (automatic),78.5,5602.25,0,66,22,32.37,6072,0,Lytle Creek,0,0,Fiber Optic,34.238162,-117.534306,1,78.5,0,4,Offer A,1090,0,0,1,0,72,1,1232.0,2330.64,0.0,5602.25,0,0,92358
5420,1,0,1,0,70,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),114.3,8244.3,0,23,30,21.68,4280,0,Mentone,1,1,Cable,34.103578000000006,-117.04054,1,114.3,0,10,Offer A,7324,1,0,1,1,70,4,0.0,1517.6,0.0,8244.3,1,1,92359
5421,0,0,0,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.05,741.5,0,33,0,41.63,2295,0,Needles,0,0,NA,34.711224,-114.702256,0,20.05,0,0,Offer C,5488,0,0,0,0,38,0,0.0,1581.94,0.0,741.5,0,0,92363
5422,1,0,1,1,68,1,0,DSL,1,1,0,0,Two year,0,Credit card (automatic),62.65,4375.8,0,38,24,36.51,5215,0,Nipton,1,1,Fiber Optic,35.478736,-115.51698400000001,1,62.65,1,4,Offer A,162,1,0,1,0,68,2,1050.0,2482.68,0.0,4375.8,0,0,92364
5423,1,0,0,0,13,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.85,1008.7,1,40,22,12.54,5964,1,San Diego,0,1,Cable,32.886925,-117.152162,0,84.084,0,0,None,74232,0,3,0,1,13,1,222.0,163.01999999999995,0.0,1008.7,0,0,92126
5424,1,1,1,0,65,1,1,Fiber optic,1,1,1,0,Two year,1,Credit card (automatic),92.7,5968.4,0,71,26,27.14,5205,0,Oro Grande,0,1,DSL,34.647959,-117.296957,1,92.7,0,3,Offer B,909,0,0,1,0,65,1,0.0,1764.1,0.0,5968.4,0,1,92368
5425,0,0,0,0,30,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,100.45,3096.9,0,27,59,34.49,3936,0,Phelan,1,0,Fiber Optic,34.441123,-117.53788600000001,0,100.45,0,0,Offer C,12463,0,0,0,1,30,1,0.0,1034.7,0.0,3096.9,1,1,92371
5426,1,0,1,0,51,1,1,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),75.2,3901.25,0,39,5,9.99,4708,0,Pinon Hills,0,1,Fiber Optic,34.459322,-117.629729,1,75.2,0,10,Offer B,4280,1,0,1,1,51,0,195.0,509.49,0.0,3901.25,0,0,92372
5427,0,0,0,0,31,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),84.75,2613.4,0,30,48,24.21,3727,0,Redlands,1,0,DSL,34.003243,-117.13828600000001,0,84.75,0,0,Offer C,31230,0,0,0,0,31,1,0.0,750.51,0.0,2613.4,0,1,92373
5428,0,0,1,0,9,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,89.45,853.1,1,62,20,26.51,4971,1,San Diego,0,0,Cable,32.886925,-117.152162,1,93.02799999999999,0,3,Offer E,74232,0,0,1,1,9,3,0.0,238.59,0.0,853.1,0,1,92126
5429,0,0,1,1,72,1,1,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),79.5,5661.7,0,35,14,32.59,4390,0,Rialto,1,0,Fiber Optic,34.109775,-117.378904,1,79.5,1,5,Offer A,75882,1,0,1,1,72,0,793.0,2346.4800000000005,0.0,5661.7,0,0,92376
5430,1,0,0,0,10,1,1,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),72.15,794.25,1,49,12,33.75,2457,1,Rialto,0,1,Fiber Optic,34.156758,-117.40468600000001,0,75.03600000000002,0,0,None,18518,0,0,0,1,10,4,95.0,337.5,0.0,794.25,0,0,92377
5431,0,0,0,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,19.8,695.05,0,62,0,30.17,5987,0,Running Springs,0,0,NA,34.186211,-117.07683,0,19.8,0,0,Offer C,5395,0,0,0,0,37,0,0.0,1116.29,0.0,695.05,0,0,92382
5432,0,0,0,0,2,1,0,DSL,0,0,1,1,Month-to-month,0,Electronic check,76.4,160.8,1,39,28,41.64,3005,1,Shoshone,1,0,Cable,35.924252,-116.18866799999999,0,79.456,0,0,Offer E,87,1,1,0,1,2,2,45.0,83.28,0.0,160.8,0,0,92384
5433,1,0,0,0,55,1,0,Fiber optic,1,1,1,1,One year,1,Mailed check,100.9,5552.05,0,19,51,42.19,5101,0,Sugarloaf,0,1,Fiber Optic,34.243088,-116.83001499999999,0,100.9,0,0,Offer B,1834,0,0,0,1,55,0,2832.0,2320.45,0.0,5552.05,1,0,92386
5434,1,0,0,1,33,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Bank transfer (automatic),95.3,3275.15,0,55,53,10.36,3087,0,Fallbrook,1,1,DSL,33.362575,-117.299644,0,95.3,3,0,Offer C,42239,0,0,0,1,33,0,0.0,341.88,0.0,3275.15,0,1,92028
5435,0,0,1,1,46,1,0,Fiber optic,0,0,0,1,One year,0,Bank transfer (automatic),90.95,4236.6,0,23,48,6.26,5187,0,Victorville,1,0,Fiber Optic,34.486835,-117.362274,1,90.95,3,2,Offer B,63235,1,0,1,1,46,1,0.0,287.96,0.0,4236.6,1,1,92392
5436,0,0,0,1,1,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,54.5,54.5,0,63,75,33.21,4359,0,Victorville,0,0,Fiber Optic,34.567058,-117.362329,0,54.5,3,0,None,12083,1,0,0,0,1,0,0.0,33.21,0.0,54.5,0,0,92394
5437,0,1,0,0,20,1,1,DSL,0,0,0,1,Month-to-month,1,Mailed check,61.6,1174.35,1,67,30,27.11,3866,1,Wrightwood,0,0,DSL,34.358321000000004,-117.61826299999998,0,64.06400000000001,0,0,None,4253,0,0,0,0,20,0,352.0,542.2,0.0,1174.35,0,0,92397
5438,1,0,1,0,9,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.9,741.7,1,35,30,19.18,4748,1,Yermo,1,1,Fiber Optic,35.013298999999996,-116.834092,1,83.096,0,0,Offer E,1195,0,1,0,0,9,7,223.0,172.62,0.0,741.7,0,0,92398
5439,1,1,0,0,32,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),96.15,3019.25,1,67,20,25.45,2246,1,Yucaipa,0,1,DSL,34.045970000000004,-117.011825,0,99.996,0,0,Offer C,41575,0,0,0,0,32,2,604.0,814.4,0.0,3019.25,0,0,92399
5440,0,0,1,1,19,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),49.6,962.9,0,43,17,7.42,5735,0,San Bernardino,1,0,Fiber Optic,34.105934999999995,-117.2914,1,49.6,1,3,None,1779,0,0,1,0,19,3,164.0,140.98,0.0,962.9,0,0,92401
5441,0,0,1,0,70,1,1,DSL,1,0,0,0,Two year,0,Credit card (automatic),65.3,4759.75,1,57,26,42.67,5591,1,San Bernardino,1,0,Cable,34.183285999999995,-117.221722,1,67.91199999999999,0,1,Offer A,53636,1,1,1,0,70,7,1238.0,2986.9,0.0,4759.75,0,0,92404
5442,0,0,0,1,61,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.0,1498.35,0,62,0,32.05,4673,0,San Bernardino,0,0,NA,34.142747,-117.30086399999999,0,25.0,1,0,Offer B,24644,0,0,0,0,61,0,0.0,1955.05,0.0,1498.35,0,0,92405
5443,1,0,0,0,26,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.45,1233.15,0,28,42,29.07,5451,0,San Bernardino,0,1,Cable,34.250069,-117.39394899999999,0,45.45,0,0,Offer C,49355,0,0,0,0,26,1,0.0,755.82,0.0,1233.15,1,1,92407
5444,1,0,1,0,45,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),107.75,4882.8,0,50,27,29.81,3301,0,San Bernardino,1,1,DSL,34.084909,-117.25810700000001,1,107.75,0,0,Offer B,12149,0,1,0,1,45,2,0.0,1341.45,0.0,4882.8,0,1,92408
5445,1,0,1,1,62,1,1,Fiber optic,0,0,1,0,Two year,1,Credit card (automatic),89.1,5411.65,0,23,73,37.75,5995,0,San Bernardino,1,1,DSL,34.106922,-117.29755300000001,1,89.1,2,4,Offer B,44556,0,0,1,0,62,0,0.0,2340.5,0.0,5411.65,1,1,92410
5446,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,19.65,1,43,0,17.25,5717,1,San Bernardino,0,1,NA,34.122501,-117.32013799999999,0,19.65,0,0,Offer E,23146,0,1,0,0,1,3,0.0,17.25,0.0,19.65,0,0,92411
5447,0,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,44.75,148.05,0,37,13,34.89,3422,0,Riverside,0,0,Fiber Optic,33.994676,-117.372498,0,44.75,0,0,None,18999,0,0,0,0,3,0,0.0,104.67,0.0,148.05,0,1,92501
5448,0,0,1,1,41,1,1,Fiber optic,1,1,0,1,One year,1,Bank transfer (automatic),101.6,3930.55,0,21,82,14.73,3275,0,Riverside,1,0,DSL,33.890046000000005,-117.455583,1,101.6,1,7,Offer B,71678,0,0,1,1,41,1,0.0,603.9300000000002,0.0,3930.55,1,1,92503
5449,1,0,1,1,67,1,0,Fiber optic,0,1,1,1,Two year,0,Bank transfer (automatic),103.15,6895.5,0,31,76,13.26,4376,0,Riverside,1,1,Cable,33.9108,-117.39815300000001,1,103.15,3,4,Offer A,46550,1,0,1,1,67,3,0.0,888.42,0.0,6895.5,0,1,92504
5450,1,0,0,0,1,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,84.65,84.65,1,25,56,22.3,4261,1,Riverside,0,1,Cable,33.920907,-117.489426,0,88.03600000000002,0,0,None,38446,0,0,0,0,1,2,0.0,22.3,0.0,84.65,1,0,92505
5451,0,0,1,0,71,1,1,Fiber optic,1,1,1,0,One year,0,Mailed check,95.65,6856.95,0,53,10,5.22,5856,0,Riverside,0,0,Fiber Optic,33.930931,-117.36178799999999,1,95.65,0,6,Offer A,42425,0,0,1,0,71,1,686.0,370.62,0.0,6856.95,0,0,92506
5452,0,0,1,1,37,1,0,DSL,1,1,1,1,One year,0,Bank transfer (automatic),75.1,2658.8,0,32,23,1.12,4131,0,Riverside,0,0,DSL,33.976328,-117.31978600000001,1,75.1,2,3,Offer C,48649,0,0,1,1,37,0,61.15,41.44000000000001,0.0,2658.8,0,1,92507
5453,1,0,1,0,60,1,0,DSL,1,1,0,0,Two year,1,Mailed check,61.35,3766.2,0,45,16,22.22,6174,0,Riverside,0,1,Cable,33.885498999999996,-117.324959,1,61.35,0,5,None,17147,1,0,1,0,60,2,603.0,1333.1999999999996,0.0,3766.2,0,0,92508
5454,0,1,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.55,69.55,1,76,24,12.46,5948,1,Riverside,0,0,Cable,34.004379,-117.447864,1,72.332,0,1,None,63999,0,6,1,0,1,3,0.0,12.46,0.0,69.55,0,0,92509
5455,0,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.7,129.55,0,50,0,31.02,5387,0,March Air Reserve Base,0,0,NA,33.888323,-117.277533,0,19.7,0,0,Offer E,1005,0,0,0,0,6,1,0.0,186.12,0.0,129.55,0,0,92518
5456,0,0,0,0,13,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,31.05,347.25,1,46,18,0.0,5131,1,Lake Elsinore,0,0,Cable,33.655421000000004,-117.391751,0,32.292,0,0,None,38519,0,2,0,0,13,4,0.0,0.0,0.0,347.25,0,1,92530
5457,0,0,1,1,11,1,0,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),51.0,581.7,0,42,57,44.84,5777,0,Lake Elsinore,0,0,Fiber Optic,33.705836,-117.31820400000001,1,51.0,3,8,None,4546,0,0,1,0,11,1,0.0,493.24,0.0,581.7,0,1,92532
5458,1,0,0,0,7,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,51.0,354.05,1,56,24,34.49,3736,1,Aguanga,0,1,Cable,33.482243,-116.827173,0,53.04,0,0,None,2433,0,0,0,0,7,2,85.0,241.43,0.0,354.05,0,0,92536
5459,0,0,1,1,10,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,88.85,929.45,0,45,51,32.76,4531,0,Anza,0,0,Fiber Optic,33.527605,-116.666551,1,88.85,3,8,None,3745,0,0,1,1,10,1,0.0,327.6,0.0,929.45,0,1,92539
5460,1,0,1,0,34,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.05,679,0,44,0,4.42,2236,0,Hemet,0,1,NA,33.739415,-116.96833899999999,1,20.05,0,6,Offer C,29687,0,0,1,0,34,2,0.0,150.28,0.0,679.0,0,0,92543
5461,0,0,0,0,62,1,0,DSL,1,0,0,1,Two year,1,Mailed check,65.1,3846.75,0,45,18,23.18,5172,0,Hemet,0,0,DSL,33.644585,-116.871544,0,65.1,0,0,None,39264,1,0,0,1,62,0,0.0,1437.16,0.0,3846.75,0,1,92544
5462,1,0,1,0,64,1,1,DSL,0,1,0,1,One year,1,Mailed check,70.15,4480.7,0,24,26,32.93,5037,0,Hemet,0,1,Fiber Optic,33.734933000000005,-117.044145,1,70.15,0,5,None,25694,1,0,1,1,64,0,0.0,2107.52,0.0,4480.7,1,1,92545
5463,0,0,1,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),44.35,44.35,1,27,65,40.42,4599,1,Homeland,0,0,Cable,33.761894,-117.12086799999999,1,46.123999999999995,3,0,None,4283,0,0,0,0,1,1,0.0,40.42,0.0,44.35,1,0,92548
5464,1,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.75,499.4,0,29,0,29.38,5161,0,Idyllwild,0,1,NA,33.755039000000004,-116.741796,0,20.75,0,0,Offer C,3588,0,1,0,0,25,2,0.0,734.5,0.0,499.4,1,0,92549
5465,0,0,0,0,26,1,0,DSL,0,1,0,0,One year,1,Mailed check,56.05,1553.2,0,30,71,35.75,3079,0,Moreno Valley,1,0,Fiber Optic,33.882740000000005,-117.224878,0,56.05,0,0,Offer C,22983,0,0,0,0,26,0,1103.0,929.5,0.0,1553.2,0,0,92551
5466,1,0,0,1,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.95,219.5,0,22,0,7.86,3044,0,Moreno Valley,0,1,NA,33.923149,-117.244933,0,19.95,1,0,None,61205,0,0,0,0,10,4,0.0,78.60000000000002,0.0,219.5,1,0,92553
5467,0,0,0,0,53,1,1,Fiber optic,1,1,1,0,One year,0,Mailed check,98.6,5311.85,0,52,12,29.39,4635,0,Moreno Valley,1,0,Fiber Optic,33.907361,-117.109972,0,98.6,0,0,None,12743,0,0,0,0,53,1,63.74,1557.67,0.0,5311.85,0,1,92555
5468,0,0,0,0,7,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.7,586.05,1,31,18,28.92,3109,1,Moreno Valley,0,0,Fiber Optic,33.970661,-117.255039,0,82.88799999999999,0,0,None,46214,0,0,0,0,7,3,105.0,202.44,0.0,586.05,0,0,92557
5469,1,0,0,0,33,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),79.0,2576.8,0,59,19,17.63,4396,0,Mountain Center,1,1,DSL,33.638645000000004,-116.55783000000001,0,79.0,0,0,Offer C,1500,0,0,0,0,33,0,0.0,581.79,0.0,2576.8,0,1,92561
5470,0,1,1,0,71,1,0,Fiber optic,0,1,0,1,Two year,0,Credit card (automatic),89.45,6435.25,0,74,27,16.26,6004,0,Murrieta,1,0,Cable,33.548869,-117.33416499999998,1,89.45,0,10,Offer A,36149,0,0,1,0,71,0,1738.0,1154.46,0.0,6435.25,0,0,92562
5471,0,0,0,0,29,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.2,1993.25,0,25,82,16.38,3982,0,Murrieta,0,0,Cable,33.581045,-117.14719,0,74.2,0,0,Offer C,18311,0,1,0,0,29,2,0.0,475.02,0.0,1993.25,1,1,92563
5472,1,0,1,1,24,1,1,DSL,1,0,1,1,Month-to-month,0,Bank transfer (automatic),81.0,1923.85,0,51,26,45.68,3019,0,Nuevo,0,1,DSL,33.827690000000004,-117.102244,1,81.0,3,3,Offer C,7344,1,0,1,1,24,0,0.0,1096.32,0.0,1923.85,0,1,92567
5473,1,0,1,1,20,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.6,939.8,0,63,10,13.18,3235,0,Perris,1,1,Fiber Optic,33.787298,-117.320676,1,49.6,1,5,None,36817,0,0,1,0,20,1,0.0,263.6,0.0,939.8,0,1,92570
5474,0,0,0,0,1,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.6,84.6,0,44,11,7.34,2196,0,Perris,0,0,Cable,33.828289,-117.20166599999999,0,84.6,0,0,Offer E,26357,0,0,0,0,1,0,0.0,7.34,0.0,84.6,0,0,92571
5475,1,0,0,1,54,1,1,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),55.0,3092.65,1,43,18,6.7,5282,1,San Jacinto,0,1,Cable,33.806708,-117.02006999999999,0,57.2,2,0,None,4456,0,0,0,0,54,3,557.0,361.8,0.0,3092.65,0,0,92582
5476,0,1,0,0,5,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,84.85,415.55,1,66,30,27.35,3305,1,San Jacinto,1,0,Fiber Optic,33.796568,-116.924723,0,88.244,0,0,None,21349,0,1,0,0,5,4,125.0,136.75,0.0,415.55,0,0,92583
5477,0,0,1,1,72,1,1,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),84.2,5986.55,0,45,53,37.84,5598,0,Menifee,1,0,DSL,33.653338,-117.178271,1,84.2,3,10,Offer A,14068,1,2,1,1,72,2,0.0,2724.4800000000005,0.0,5986.55,0,1,92584
5478,1,0,1,0,52,1,0,Fiber optic,1,1,1,1,Two year,1,Electronic check,106.3,5487,0,26,51,49.82,4969,0,Sun City,1,1,Fiber Optic,33.739412,-117.17333400000001,1,106.3,0,4,None,8692,1,0,1,1,52,0,0.0,2590.64,0.0,5487.0,1,1,92585
5479,0,0,0,0,9,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.05,651.5,0,63,5,29.87,5121,0,Sun City,0,0,Fiber Optic,33.707483,-117.200006,0,69.05,0,0,Offer E,18161,0,0,0,0,9,0,0.0,268.83,0.0,651.5,0,1,92586
5480,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.4,45.4,0,38,21,49.33,4916,0,Sun City,0,0,Fiber Optic,33.69887,-117.25071000000001,0,45.4,0,0,Offer E,13151,0,0,0,0,1,0,0.0,49.33,0.0,45.4,0,0,92587
5481,1,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.65,73.65,1,80,21,39.88,5443,1,Temecula,0,1,Cable,33.475493,-117.219551,0,76.596,0,0,None,3070,0,0,0,0,1,4,0.0,39.88,0.0,73.65,0,0,92590
5482,1,0,1,1,33,1,0,DSL,0,0,1,1,One year,1,Mailed check,73.9,2405.05,1,33,4,33.32,5374,1,Temecula,1,1,Cable,33.540603999999995,-117.10909,1,76.85600000000002,0,3,Offer C,25655,1,1,1,1,33,3,96.0,1099.56,0.0,2405.05,0,0,92591
5483,0,0,1,0,55,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,77.75,4458.15,1,38,4,19.41,4398,1,Temecula,1,0,Cable,33.507255,-117.029473,1,80.86,0,5,None,46171,0,1,1,0,55,1,178.0,1067.55,0.0,4458.15,0,0,92592
5484,1,0,1,1,69,1,1,Fiber optic,0,0,1,1,Two year,1,Electronic check,99.35,6856.45,0,55,21,8.46,4637,0,Wildomar,0,1,Cable,33.617108,-117.253349,1,99.35,1,0,Offer A,19368,1,0,0,1,69,0,1440.0,583.74,0.0,6856.45,0,0,92595
5485,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,50.75,50.75,0,37,20,45.77,2250,0,Winchester,0,1,Fiber Optic,33.657433000000005,-117.04253999999999,0,50.75,0,0,Offer E,4093,0,0,0,0,1,1,0.0,45.77,0.0,50.75,0,1,92596
5486,1,0,0,0,54,1,1,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),87.1,4735.2,0,60,26,18.54,5418,0,Irvine,1,1,Cable,33.720359,-117.733655,0,87.1,0,0,None,2762,1,0,0,1,54,2,1231.0,1001.16,0.0,4735.2,0,0,92602
5487,1,0,0,1,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.15,682.15,0,51,0,21.16,5759,0,Irvine,0,1,NA,33.688546,-117.788091,0,20.15,3,0,Offer C,27369,0,0,0,0,33,1,0.0,698.28,0.0,682.15,0,0,92604
5488,1,1,1,0,45,1,1,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),98.7,4525.8,0,71,20,2.38,2535,0,Irvine,1,1,Fiber Optic,33.703976000000004,-117.82417199999999,1,98.7,0,1,Offer B,17621,1,1,1,0,45,1,0.0,107.1,0.0,4525.8,0,1,92606
5489,0,0,0,1,11,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,25.2,321.05,0,49,19,0.0,5916,0,Foothill Ranch,0,0,Fiber Optic,33.698728,-117.67768000000001,0,25.2,1,0,None,10936,0,0,0,0,11,0,0.0,0.0,0.0,321.05,0,1,92610
5490,1,0,0,0,6,1,0,DSL,1,1,0,0,Month-to-month,1,Bank transfer (automatic),55.7,335.65,0,22,41,3.16,2482,0,Irvine,0,1,Fiber Optic,33.643095,-117.810896,0,55.7,0,0,None,41062,0,0,0,0,6,0,13.76,18.96,0.0,335.65,1,1,92612
5491,1,0,0,0,21,1,0,DSL,1,0,1,0,Month-to-month,0,Bank transfer (automatic),65.35,1424.4,0,28,42,16.16,2887,0,Irvine,1,1,Fiber Optic,33.680302000000005,-117.83329599999999,0,65.35,0,0,None,22499,0,0,0,0,21,0,0.0,339.36,0.0,1424.4,1,1,92614
5492,0,0,1,1,65,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.3,1748.55,0,25,0,34.03,4533,0,Irvine,0,0,NA,33.667145,-117.73213500000001,1,25.3,3,9,None,6301,0,0,1,0,65,1,0.0,2211.9500000000007,0.0,1748.55,1,0,92618
5493,0,1,1,0,6,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.35,474.9,1,78,19,28.71,5721,1,Irvine,0,0,DSL,33.716136,-117.752574,1,87.72399999999999,0,1,None,26419,0,0,1,0,6,0,90.0,172.26,0.0,474.9,0,0,92620
5494,0,0,0,0,8,1,0,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,84.95,668.4,1,35,7,32.31,4437,1,Capistrano Beach,0,0,Fiber Optic,33.458754,-117.665104,0,88.348,0,0,None,7465,0,0,0,0,8,3,47.0,258.48,0.0,668.4,0,0,92624
5495,1,0,0,0,11,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.85,926.25,1,40,28,44.94,3634,1,Corona Del Mar,0,1,Fiber Optic,33.600986999999996,-117.862734,0,76.804,0,0,None,13422,1,2,0,0,11,4,259.0,494.34,0.0,926.25,0,0,92625
5496,1,0,1,1,43,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.25,1077.95,0,60,0,2.81,4432,0,Costa Mesa,0,1,NA,33.678591,-117.90547099999999,1,24.25,2,4,None,48207,0,0,1,0,43,0,0.0,120.83,0.0,1077.95,0,0,92626
5497,1,0,1,1,49,0,No phone service,DSL,0,1,1,1,One year,1,Bank transfer (automatic),51.8,2541.25,1,57,6,0.0,5375,1,Costa Mesa,0,1,Cable,33.645672,-117.92261299999998,1,53.872,0,2,None,62069,0,1,1,1,49,4,152.0,0.0,0.0,2541.25,0,0,92627
5498,0,1,1,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,46.0,46,1,69,21,7.74,4531,1,Dana Point,0,0,Cable,33.477923,-117.70531399999999,1,47.84,0,1,None,27730,0,0,1,0,1,0,0.0,7.74,0.0,46.0,0,0,92629
5499,1,1,0,0,15,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.4,1156.1,1,78,13,17.23,3621,1,Lake Forest,0,1,DSL,33.644849,-117.68425400000001,0,82.57600000000002,0,0,None,59176,0,0,0,0,15,0,150.0,258.45,0.0,1156.1,0,0,92630
5500,1,0,1,1,60,1,0,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),60.5,3694.45,0,37,28,43.24,6026,0,Huntington Beach,1,1,DSL,33.666301000000004,-117.969501,1,60.5,2,7,None,56517,0,0,1,0,60,1,1034.0,2594.4,0.0,3694.45,0,0,92646
5501,1,0,0,0,17,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),25.1,382.8,0,48,11,0.0,4580,0,Huntington Beach,0,1,DSL,33.723579,-118.00544099999999,0,25.1,0,0,None,58764,0,1,0,0,17,1,42.0,0.0,0.0,382.8,0,0,92647
5502,1,1,1,0,16,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),71.8,1167.8,1,78,6,45.9,3327,1,Huntington Beach,0,1,Cable,33.679659,-118.016195,1,74.672,0,1,None,42663,0,0,1,0,16,0,70.0,734.4,0.0,1167.8,0,0,92648
5503,1,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.05,746.75,0,24,0,41.02,3942,0,Huntington Beach,0,1,NA,33.721917,-118.043237,1,20.05,1,4,Offer C,32304,0,0,1,0,35,1,0.0,1435.7,0.0,746.75,1,0,92649
5504,1,1,1,0,44,1,1,Fiber optic,0,1,0,1,One year,0,Mailed check,88.4,3912.9,1,68,15,24.62,2674,1,Laguna Beach,0,1,DSL,33.570023,-117.773669,1,91.936,0,1,None,25206,0,0,1,1,44,0,587.0,1083.28,0.0,3912.9,0,0,92651
5505,0,0,1,1,12,0,No phone service,DSL,0,0,0,0,One year,0,Credit card (automatic),30.25,368.85,0,48,22,0.0,5988,0,Laguna Hills,0,0,Cable,33.606899,-117.717854,1,30.25,1,4,None,48273,1,1,1,0,12,2,81.0,0.0,0.0,368.85,0,0,92653
5506,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.2,20.2,0,63,0,13.08,4496,0,Midway City,0,1,NA,33.744439,-117.98588000000001,0,20.2,0,0,None,8660,0,0,0,0,1,0,0.0,13.08,0.0,20.2,0,0,92655
5507,0,0,0,0,28,1,0,DSL,1,1,0,0,One year,1,Electronic check,59.9,1654.7,0,57,11,11.32,4131,0,Aliso Viejo,0,0,DSL,33.571259000000005,-117.731917,0,59.9,0,0,Offer C,41237,1,0,0,0,28,0,0.0,316.9600000000001,0.0,1654.7,0,1,92656
5508,1,0,1,0,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.15,1940.85,0,61,0,9.03,4279,0,Newport Coast,0,1,NA,33.603282,-117.82184099999999,1,25.15,0,7,Offer A,5597,0,0,1,0,70,0,0.0,632.0999999999998,0.0,1940.85,0,0,92657
5509,0,0,0,1,5,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,46.0,221.7,1,56,15,23.89,4846,1,Newport Beach,0,0,Cable,33.634626000000004,-117.874882,0,47.84,1,0,None,28687,0,0,0,0,5,0,33.0,119.45,0.0,221.7,0,0,92660
5510,1,0,0,0,18,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Credit card (automatic),101.3,1794.65,0,61,20,7.56,5948,0,Newport Beach,1,1,Fiber Optic,33.601309,-117.902304,0,101.3,0,0,None,4242,0,0,0,1,18,1,0.0,136.07999999999998,0.0,1794.65,0,1,92661
5511,1,0,1,0,70,1,1,DSL,1,0,1,1,Two year,1,Credit card (automatic),76.95,5289.8,0,46,18,18.26,6280,0,Newport Beach,0,1,DSL,33.606336,-117.893042,1,76.95,0,1,Offer A,3124,1,0,1,1,70,0,95.22,1278.2,0.0,5289.8,0,1,92662
5512,0,0,1,1,9,1,1,DSL,0,1,0,0,Month-to-month,1,Mailed check,55.3,501.2,0,51,22,23.36,4291,0,Newport Beach,0,0,Fiber Optic,33.62251,-117.927024,1,55.3,3,1,None,22133,0,0,1,0,9,0,0.0,210.24,0.0,501.2,0,1,92663
5513,0,1,0,0,67,1,0,Fiber optic,1,1,1,0,Two year,1,Bank transfer (automatic),92.45,6140.85,0,69,21,2.57,5857,0,San Clemente,0,0,Fiber Optic,33.429488,-117.60943200000001,0,92.45,0,0,Offer A,34946,1,0,0,0,67,0,0.0,172.19,0.0,6140.85,0,1,92672
5514,0,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),48.45,48.45,0,63,21,16.42,5838,0,San Clemente,0,0,Fiber Optic,33.4725,-117.584273,0,48.45,0,0,None,15297,0,1,0,0,1,1,0.0,16.42,0.0,48.45,0,1,92673
5515,0,0,1,1,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.35,309.25,0,20,0,20.0,2269,0,San Juan Capistrano,0,0,NA,33.521446999999995,-117.60255500000001,1,19.35,3,5,None,34321,0,0,1,0,18,0,0.0,360.0,0.0,309.25,1,0,92675
5516,1,0,0,0,4,1,1,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),51.75,201.1,1,39,14,9.98,3865,1,Silverado,0,1,DSL,33.782346000000004,-117.635263,0,53.82,0,0,None,1859,0,2,0,0,4,1,28.0,39.92,0.0,201.1,0,0,92676
5517,1,1,1,1,71,1,0,Fiber optic,1,1,0,0,One year,1,Bank transfer (automatic),86.7,6179.35,0,76,19,30.16,4485,0,Laguna Niguel,1,1,DSL,33.529047,-117.701175,1,86.7,2,5,Offer A,62103,0,0,1,0,71,0,1174.0,2141.36,0.0,6179.35,0,0,92677
5518,1,0,1,1,30,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,94.4,2838.7,1,52,7,28.85,2792,1,Trabuco Canyon,0,1,DSL,33.631119,-117.567346,1,98.17600000000002,0,1,Offer C,32268,0,0,1,0,30,3,199.0,865.5,0.0,2838.7,0,0,92679
5519,1,0,1,0,1,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,55.7,55.7,0,61,9,17.68,5664,0,Westminster,1,1,DSL,33.752590999999995,-117.99366100000002,1,55.7,0,10,None,88230,0,0,1,0,1,1,0.0,17.68,0.0,55.7,0,0,92683
5520,0,0,0,0,55,1,1,Fiber optic,1,0,0,0,One year,1,Credit card (automatic),84.25,4589.85,0,19,48,44.85,5735,0,Rancho Santa Margarita,1,0,DSL,33.624654,-117.611733,0,84.25,0,0,None,42193,0,0,0,0,55,0,2203.0,2466.75,0.0,4589.85,1,0,92688
5521,1,0,0,0,59,1,0,DSL,0,0,1,0,Month-to-month,1,Electronic check,64.65,3735.45,0,60,18,16.8,5687,0,Mission Viejo,1,1,Cable,33.611945,-117.66586699999999,0,64.65,0,0,None,46371,1,0,0,0,59,0,0.0,991.2,0.0,3735.45,0,1,92691
5522,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.15,70.15,1,34,7,2.24,3208,1,Mission Viejo,0,0,Cable,33.60693,-117.644253,0,72.956,0,0,None,46227,0,0,0,0,1,0,0.0,2.24,0.0,70.15,0,0,92692
5523,0,0,1,0,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.2,477.55,0,19,73,41.22,2551,0,Ladera Ranch,0,0,Fiber Optic,33.569186,-117.640055,1,69.2,0,8,None,350,0,0,1,0,7,2,0.0,288.54,0.0,477.55,1,1,92694
5524,1,0,1,1,45,1,0,DSL,1,0,0,0,Two year,0,Bank transfer (automatic),54.65,2553.7,0,21,59,45.21,5083,0,Santa Ana,0,1,DSL,33.748478000000006,-117.85891799999999,1,54.65,1,1,None,58157,1,0,1,0,45,0,150.67,2034.45,0.0,2553.7,1,1,92701
5525,0,0,1,1,54,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),24.75,1342.15,0,40,0,28.87,6466,0,Santa Ana,0,0,NA,33.748635,-117.906125,1,24.75,2,1,None,70011,0,0,1,0,54,2,0.0,1558.98,0.0,1342.15,0,0,92703
5526,1,0,1,1,51,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,23.95,1216.35,0,40,0,42.55,5895,0,Santa Ana,0,1,NA,33.719869,-117.907063,1,23.95,3,1,None,91188,0,0,1,0,51,0,0.0,2170.05,0.0,1216.35,0,0,92704
5527,0,1,1,0,72,1,1,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),105.0,7578.05,0,78,10,27.79,6423,0,Santa Ana,1,0,Fiber Optic,33.766003999999995,-117.786763,1,105.0,0,1,Offer A,44117,0,0,1,0,72,1,758.0,2000.88,0.0,7578.05,0,0,92705
5528,1,0,1,0,44,1,0,DSL,1,1,0,0,One year,1,Bank transfer (automatic),59.85,2603.95,0,39,24,17.61,5981,0,Santa Ana,0,1,Fiber Optic,33.765893,-117.881533,1,59.85,0,1,None,37879,1,0,1,0,44,0,625.0,774.8399999999998,0.0,2603.95,0,0,92706
5529,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,42.7,0,19,0,40.28,4394,0,Santa Ana,0,1,NA,33.714828999999995,-117.872941,0,20.05,0,0,None,62634,0,0,0,0,2,1,0.0,80.56,0.0,42.7,1,0,92707
5530,0,0,0,0,66,1,1,Fiber optic,0,0,1,0,One year,1,Bank transfer (automatic),92.15,6056.9,0,49,28,19.68,4928,0,Fountain Valley,1,0,DSL,33.712036,-117.95011299999999,0,92.15,0,0,Offer A,54548,0,0,0,0,66,0,1696.0,1298.88,0.0,6056.9,0,0,92708
5531,1,0,1,1,68,0,No phone service,DSL,1,1,1,0,One year,0,Mailed check,44.8,2983.65,0,39,19,0.0,4112,0,Tustin,0,1,Cable,33.735802,-117.818805,1,44.8,2,1,Offer A,55062,0,0,1,0,68,1,567.0,0.0,0.0,2983.65,0,0,92780
5532,0,0,0,0,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.9,689.35,0,52,0,26.16,5581,0,Tustin,0,0,NA,33.738543,-117.785046,0,20.9,0,0,None,17494,0,0,0,0,31,0,0.0,810.96,0.0,689.35,0,0,92782
5533,0,1,0,0,21,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.4,2025.1,0,77,16,37.4,5691,0,Anaheim,0,0,Fiber Optic,33.844983,-117.952151,0,95.4,0,0,None,60553,0,1,0,0,21,1,0.0,785.4,0.0,2025.1,0,1,92801
5534,1,0,0,1,21,1,1,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,80.35,1747.2,0,61,24,13.39,4579,0,Anaheim,0,1,Cable,33.807864,-117.923782,0,80.35,2,0,Offer D,45086,0,0,0,0,21,0,419.0,281.19,0.0,1747.2,0,0,92802
5535,0,0,1,1,55,1,1,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),85.1,4657.95,0,37,52,8.39,5661,0,Anaheim,1,0,Fiber Optic,33.818000000000005,-117.974404,1,85.1,3,1,None,81333,1,1,1,1,55,2,2422.0,461.4500000000001,0.0,4657.95,0,0,92804
5536,1,0,0,0,9,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),34.7,296.1,1,43,10,0.0,5352,1,Anaheim,0,1,Cable,33.830209,-117.906099,0,36.088,0,0,None,68802,0,0,0,0,9,2,0.0,0.0,0.0,296.1,0,1,92805
5537,1,1,1,0,71,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),115.05,8016.6,0,72,18,46.82,4438,0,Anaheim,1,1,Fiber Optic,33.837959999999995,-117.870494,1,115.05,0,1,Offer A,34398,1,0,1,0,71,0,0.0,3324.22,0.0,8016.6,0,1,92806
5538,0,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,81.1,81.1,1,53,26,22.86,2075,1,Anaheim,0,0,Fiber Optic,33.848733,-117.788357,0,84.344,0,0,None,36301,0,0,0,1,1,2,0.0,22.86,0.0,81.1,0,0,92807
5539,1,0,1,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.95,433.5,0,37,0,37.4,2233,0,Anaheim,0,1,NA,33.850452000000004,-117.72666799999999,1,19.95,1,1,Offer D,19629,0,0,1,0,22,2,0.0,822.8,0.0,433.5,0,0,92808
5540,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.55,20.55,1,25,0,37.92,3797,1,Brea,0,0,NA,33.930199,-117.862898,1,20.55,2,1,None,34055,0,0,1,0,1,1,0.0,37.92,0.0,20.55,1,0,92821
5541,0,0,0,0,61,1,1,Fiber optic,0,0,1,1,Two year,1,Electronic check,106.6,6428.4,1,39,31,41.23,4183,1,Brea,1,0,Cable,33.924143,-117.79387,0,110.86399999999999,0,0,None,1408,1,1,0,1,61,2,1993.0,2515.03,0.0,6428.4,0,0,92823
5542,0,0,1,0,67,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),86.15,5883.85,0,41,23,3.2,5037,0,Fullerton,1,0,DSL,33.879983,-117.895482,1,86.15,0,1,Offer A,34592,1,1,1,1,67,1,135.33,214.4,0.0,5883.85,0,1,92831
5543,0,1,0,0,14,1,0,Fiber optic,1,1,0,0,Month-to-month,0,Electronic check,78.85,1043.8,0,76,2,48.01,5327,0,Fullerton,0,0,Cable,33.868316,-117.929029,0,78.85,0,0,None,24502,0,0,0,0,14,1,0.0,672.14,0.0,1043.8,0,1,92832
5544,1,0,1,0,59,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,106.75,6252.9,1,47,23,49.31,4508,1,Fullerton,1,1,Cable,33.877639,-117.96121200000002,1,111.02,0,7,None,46105,1,1,1,0,59,3,1438.0,2909.29,0.0,6252.9,0,0,92833
5545,1,1,1,0,21,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Bank transfer (automatic),86.55,1857.25,0,71,9,22.3,5318,0,Fullerton,1,1,Fiber Optic,33.902211,-117.914922,1,86.55,0,0,None,21157,0,0,0,0,21,1,0.0,468.3,0.0,1857.25,0,1,92835
5546,1,0,0,0,4,0,No phone service,DSL,1,1,0,0,Month-to-month,0,Mailed check,42.4,146.4,0,50,23,0.0,4282,0,Garden Grove,0,1,DSL,33.787165,-117.93188899999998,0,42.4,0,0,None,50641,1,0,0,0,4,0,3.37,0.0,0.0,146.4,0,1,92840
5547,0,0,0,0,3,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.45,240.45,1,56,14,16.15,3591,1,Garden Grove,0,0,DSL,33.786738,-117.982564,0,93.02799999999999,0,0,None,31428,0,0,0,1,3,3,0.0,48.45,0.0,240.45,0,1,92841
5548,1,0,1,0,70,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.25,1724.15,0,36,0,28.54,4118,0,Garden Grove,0,1,NA,33.764018,-117.93150700000001,1,24.25,0,1,Offer A,43491,0,0,1,0,70,1,0.0,1997.8,0.0,1724.15,0,0,92843
5549,0,0,0,0,3,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,97.9,315.3,1,40,8,30.18,4330,1,Garden Grove,0,0,Cable,33.766476000000004,-117.96979499999999,0,101.816,0,0,None,23481,1,0,0,1,3,0,25.0,90.54,0.0,315.3,0,0,92844
5550,1,1,0,0,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.5,429.55,0,79,0,23.23,5766,0,Garden Grove,0,1,NA,33.782955,-118.02645600000001,0,20.5,0,0,None,15878,0,0,0,0,21,1,0.0,487.83,0.0,429.55,0,0,92845
5551,1,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.6,356.15,0,46,0,29.12,5909,0,Norco,0,1,NA,33.925833000000004,-117.55963899999999,0,19.6,0,0,Offer D,22443,0,0,0,0,20,2,0.0,582.4,0.0,356.15,0,0,92860
5552,1,0,1,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.25,488.25,0,50,0,37.7,3339,0,Villa Park,0,1,NA,33.817473,-117.81046200000002,1,20.25,2,1,Offer D,5935,0,0,1,0,22,3,0.0,829.4000000000002,0.0,488.25,0,0,92861
5553,1,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,1,Mailed check,55.7,55.7,1,62,24,48.22,4629,1,Orange,0,1,DSL,33.828779,-117.848299,0,57.928,0,0,None,18058,0,1,0,1,1,5,0.0,48.22,0.0,55.7,0,0,92865
5554,0,0,0,0,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.6,1298.7,0,25,0,16.57,6469,0,Orange,0,0,NA,33.784597,-117.84453500000001,0,20.6,0,0,None,15396,0,0,0,0,63,1,0.0,1043.91,0.0,1298.7,1,0,92866
5555,0,0,1,1,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.8,1378.75,0,38,0,48.44,5169,0,Orange,0,0,NA,33.81859,-117.821288,1,19.8,2,1,Offer A,40915,0,0,1,0,70,0,0.0,3390.8,0.0,1378.75,0,0,92867
5556,1,0,0,0,13,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.8,973.45,1,61,3,30.88,5067,1,Orange,1,1,Cable,33.787796,-117.875928,0,82.992,0,0,None,23172,0,1,0,0,13,1,0.0,401.44,0.0,973.45,0,1,92868
5557,0,0,0,0,5,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,80.2,384.25,0,25,59,48.86,3391,0,Orange,0,0,Cable,33.792790999999994,-117.789749,0,80.2,0,0,Offer E,37916,0,0,0,0,5,2,0.0,244.3,0.0,384.25,1,1,92869
5558,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),116.4,8543.25,0,61,20,28.86,6491,0,Placentia,1,0,DSL,33.881158,-117.85478300000001,1,116.4,2,1,Offer A,48170,1,0,1,1,72,1,0.0,2077.92,0.0,8543.25,0,1,92870
5559,0,0,0,0,13,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,31.65,389.95,0,27,27,0.0,4959,0,Corona,0,0,Fiber Optic,33.893823,-117.531446,0,31.65,0,0,Offer D,44875,0,0,0,0,13,0,105.0,0.0,0.0,389.95,1,0,92879
5560,1,0,1,0,61,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Credit card (automatic),94.15,5731.85,0,63,2,17.73,4806,0,Corona,1,1,Cable,33.918043,-117.61780900000001,1,94.15,0,1,None,16998,1,0,1,1,61,1,115.0,1081.53,0.0,5731.85,0,0,92880
5561,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.65,20.65,0,50,0,1.47,2729,0,Corona,0,1,NA,33.833686,-117.51306299999999,0,20.65,0,0,Offer E,21911,0,0,0,0,1,0,0.0,1.47,0.0,20.65,0,0,92881
5562,0,1,1,0,56,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),76.85,4275.75,0,72,29,27.56,6035,0,Corona,0,0,DSL,33.819385,-117.60021299999998,1,76.85,0,7,Offer B,60294,1,0,1,0,56,2,1240.0,1543.36,0.0,4275.75,0,0,92882
5563,0,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.15,84.5,0,35,0,32.54,5535,0,Corona,0,0,NA,33.762351,-117.488725,0,20.15,0,0,Offer E,13188,0,0,0,0,4,2,0.0,130.16,0.0,84.5,0,0,92883
5564,1,0,0,0,35,1,1,DSL,1,0,0,0,Two year,0,Mailed check,55.25,1924.1,0,64,21,20.39,5498,0,Yorba Linda,0,1,Fiber Optic,33.897253000000006,-117.792202,0,55.25,0,0,None,39458,0,1,0,0,35,1,0.0,713.65,0.0,1924.1,0,1,92886
5565,0,0,1,0,18,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,39.05,669.85,1,46,33,0.0,2601,1,Yorba Linda,1,0,Fiber Optic,33.884073,-117.732197,1,40.611999999999995,0,1,None,20893,0,1,1,0,18,2,221.0,0.0,0.0,669.85,0,0,92887
5566,1,0,1,0,72,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),82.15,5784.3,0,62,5,22.01,4552,0,Ventura,1,1,DSL,34.360261,-119.30638300000001,1,82.15,0,5,Offer A,32899,0,0,1,1,72,1,28.92,1584.72,0.0,5784.3,0,1,93001
5567,0,1,0,0,49,1,1,Fiber optic,1,1,0,1,One year,0,Bank transfer (automatic),103.0,5166.2,0,77,21,36.47,5023,0,Ventura,1,0,Cable,34.279221,-119.22143700000001,0,103.0,0,0,Offer B,46894,1,0,0,1,49,4,0.0,1787.03,0.0,5166.2,0,1,93003
5568,0,0,1,0,44,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),95.1,4060.55,0,46,6,32.72,2221,0,Ventura,1,0,Cable,34.278696999999994,-119.167798,1,95.1,0,10,Offer B,27381,1,0,1,0,44,0,244.0,1439.6799999999996,0.0,4060.55,0,0,93004
5569,0,1,1,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,83.9,267.4,1,75,12,7.38,3464,1,Camarillo,0,0,Cable,34.227846,-119.079903,1,87.25600000000001,0,3,None,42853,1,3,1,0,3,1,32.0,22.14,0.0,267.4,0,0,93010
5570,0,0,1,1,37,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,95.15,3532.85,0,40,15,41.03,3407,0,Camarillo,1,0,Fiber Optic,34.205504,-118.99311100000001,1,95.15,1,2,None,24945,0,0,1,1,37,1,530.0,1518.11,0.0,3532.85,0,0,93012
5571,1,0,1,0,61,1,1,DSL,0,1,1,1,One year,1,Electronic check,79.8,4914.8,0,36,5,27.88,6432,0,Carpinteria,1,1,DSL,34.441398,-119.51316299999999,1,79.8,0,7,Offer B,17409,0,0,1,1,61,0,0.0,1700.6799999999996,0.0,4914.8,0,1,93013
5572,1,0,1,0,70,1,1,DSL,1,0,0,1,Two year,1,Credit card (automatic),74.8,5315.8,0,34,5,8.28,6447,0,Fillmore,1,1,Fiber Optic,34.408161,-118.86511100000001,1,74.8,0,9,Offer A,16013,1,0,1,1,70,0,266.0,579.5999999999998,0.0,5315.8,0,0,93015
5573,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.85,69.85,1,70,33,43.45,5056,1,Moorpark,0,0,Cable,34.312945,-118.85816899999999,0,72.64399999999998,0,0,None,32984,0,0,0,0,1,1,0.0,43.45,0.0,69.85,0,0,93021
5574,0,0,0,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.45,775.6,0,52,0,15.48,2839,0,Oak View,0,0,NA,34.404544,-119.302118,0,20.45,0,0,Offer B,6503,0,0,0,0,41,0,0.0,634.6800000000002,0.0,775.6,0,0,93022
5575,1,0,1,1,70,1,1,DSL,1,1,0,1,One year,0,Bank transfer (automatic),78.35,5445.95,0,25,59,35.9,4422,0,Ojai,1,1,Fiber Optic,34.581308,-118.93194799999999,1,78.35,1,2,Offer A,21633,1,0,1,1,70,0,0.0,2513.0,0.0,5445.95,1,1,93023
5576,0,0,0,0,1,1,0,DSL,0,0,1,0,Month-to-month,1,Mailed check,53.55,53.55,1,61,15,1.59,2326,1,Oxnard,0,0,Fiber Optic,34.223244,-119.18012,0,55.692,0,0,None,79736,0,0,0,0,1,5,0.0,1.59,0.0,53.55,0,0,93030
5577,1,0,0,0,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,19.1,1007.8,0,34,0,29.33,4120,0,Oxnard,0,1,NA,34.156628999999995,-119.117218,0,19.1,0,0,Offer B,77791,0,1,0,0,51,2,0.0,1495.83,0.0,1007.8,0,0,93033
5578,0,0,1,1,42,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.0,833.55,0,63,0,3.14,3413,0,Oxnard,0,0,NA,34.184540000000005,-119.22466599999998,1,20.0,1,3,Offer B,25322,0,1,1,0,42,2,0.0,131.88,0.0,833.55,0,0,93035
5579,0,0,1,1,70,1,1,Fiber optic,1,1,0,0,Two year,0,Bank transfer (automatic),93.9,6579.05,1,38,15,5.48,6173,1,Piru,1,0,DSL,34.432843,-118.730106,1,97.656,0,1,Offer A,1459,1,0,1,0,70,1,0.0,383.6,0.0,6579.05,0,1,93040
5580,1,0,0,0,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.95,1004.5,0,43,0,11.02,4254,0,Port Hueneme,0,1,NA,34.110124,-119.100972,0,19.95,0,0,Offer B,25634,0,1,0,0,48,3,0.0,528.96,0.0,1004.5,0,0,93041
5581,1,0,1,1,68,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,113.15,7856,1,48,24,23.67,4610,1,Santa Paula,1,1,Cable,34.402343,-119.094824,1,117.67600000000002,0,1,Offer A,32511,1,0,1,1,68,2,1885.0,1609.5600000000004,0.0,7856.0,0,0,93060
5582,0,0,0,0,48,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.0,1183.05,0,54,0,30.82,3948,0,Simi Valley,0,0,NA,34.296813,-118.685703,0,24.0,0,0,Offer B,49027,0,0,0,0,48,2,0.0,1479.36,0.0,1183.05,0,0,93063
5583,0,1,1,0,26,1,0,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,84.95,2169.75,1,65,3,18.26,4316,1,Simi Valley,0,0,DSL,34.269449,-118.76847099999999,1,88.348,0,1,Offer C,64802,0,0,1,1,26,1,0.0,474.7600000000001,0.0,2169.75,0,1,93065
5584,1,0,1,0,11,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.5,896.9,1,42,30,11.5,5119,1,Somis,0,1,Cable,34.297628,-119.014627,1,83.72,0,3,Offer D,2966,0,1,1,0,11,1,0.0,126.5,0.0,896.9,0,1,93066
5585,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.3,19.3,1,61,0,49.2,4266,1,Summerland,0,1,NA,34.420998,-119.60136999999999,0,19.3,0,0,None,576,0,4,0,0,1,1,0.0,49.2,0.0,19.3,0,0,93067
5586,0,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.15,501.35,0,36,0,20.18,5606,0,Santa Barbara,0,0,NA,34.419203,-119.710008,0,19.15,0,0,None,31727,0,0,0,0,27,1,0.0,544.86,0.0,501.35,0,0,93101
5587,0,1,0,0,46,1,0,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),91.3,4126.35,0,65,26,11.93,3191,0,Santa Barbara,1,0,Fiber Optic,34.438581,-119.685368,0,91.3,0,0,Offer B,20893,0,0,0,0,46,2,0.0,548.78,0.0,4126.35,0,1,93103
5588,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,49.65,49.65,1,60,9,4.18,5338,1,Santa Barbara,1,1,DSL,34.037341999999995,-119.80078999999999,0,51.636,0,0,None,25771,0,0,0,0,1,5,0.0,4.18,0.0,49.65,0,0,93105
5589,0,0,0,0,46,1,0,DSL,0,0,0,0,Two year,0,Credit card (automatic),54.35,2460.15,1,52,19,45.2,2793,1,Santa Barbara,1,0,DSL,34.457541,-119.631072,0,56.523999999999994,0,0,None,12741,1,5,0,0,46,3,467.0,2079.2000000000007,0.0,2460.15,0,0,93108
5590,1,0,1,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.15,477.6,0,49,0,19.09,3829,0,Santa Barbara,0,1,NA,34.406256,-119.72693600000001,1,19.15,2,5,None,10986,0,0,1,0,25,0,0.0,477.25,0.0,477.6,0,0,93109
5591,1,0,0,0,4,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,88.45,370.65,1,32,16,49.14,2456,1,Santa Barbara,0,1,DSL,34.437945,-119.77191,0,91.988,0,0,None,15757,0,1,0,1,4,2,0.0,196.56,0.0,370.65,0,1,93110
5592,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,265.75,0,56,0,10.11,2016,0,Santa Barbara,0,1,NA,34.460196999999994,-119.80260200000001,0,19.75,0,0,Offer D,16477,0,1,0,0,13,2,0.0,131.43,0.0,265.75,0,0,93111
5593,1,0,1,0,31,1,0,DSL,1,1,0,1,One year,1,Credit card (automatic),75.5,2424.45,0,41,15,27.37,5611,0,Goleta,1,1,Cable,34.489983,-120.091246,1,75.5,0,2,None,49975,1,0,1,1,31,1,36.37,848.47,0.0,2424.45,0,1,93117
5594,0,0,1,1,23,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,83.75,1849.95,0,30,30,34.91,3585,0,Alpaugh,0,0,Fiber Optic,35.869626000000004,-119.49877099999999,1,83.75,2,1,Offer D,1054,0,0,1,0,23,1,555.0,802.93,0.0,1849.95,0,0,93201
5595,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.4,61.05,0,58,0,6.65,5816,0,Armona,0,0,NA,36.315979,-119.710852,0,19.4,0,0,None,2872,0,0,0,0,2,0,0.0,13.3,0.0,61.05,0,0,93202
5596,0,0,0,0,65,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),26.5,1698.55,0,42,0,33.71,4404,0,Arvin,0,0,NA,35.116307,-118.817644,0,26.5,0,0,Offer B,16206,0,1,0,0,65,1,0.0,2191.15,0.0,1698.55,0,0,93203
5597,1,1,0,0,22,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),90.5,1910.6,1,71,30,46.11,5014,1,Avenal,0,1,Fiber Optic,35.916942999999996,-120.129921,0,94.12,0,0,None,14697,1,1,0,0,22,4,573.0,1014.42,0.0,1910.6,0,0,93204
5598,0,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.15,998.1,0,31,0,27.7,5390,0,Bodfish,0,0,NA,35.523990999999995,-118.40043200000001,1,19.15,1,0,Offer B,1954,0,0,0,0,55,0,0.0,1523.5,0.0,998.1,0,0,93205
5599,1,0,1,0,9,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Mailed check,94.85,890.6,1,54,7,17.47,3016,1,Buttonwillow,1,1,DSL,35.451402,-119.488413,1,98.644,0,1,None,2078,1,0,1,0,9,2,62.0,157.23,0.0,890.6,0,0,93206
5600,1,0,1,1,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),69.95,529.5,1,49,3,35.42,3296,1,California Hot Springs,0,1,DSL,35.865795,-118.69758999999999,1,72.748,0,9,None,226,0,0,1,0,7,4,16.0,247.94,0.0,529.5,0,0,93207
5601,0,0,1,1,35,0,No phone service,DSL,0,0,1,0,One year,0,Mailed check,40.9,1383.6,0,36,30,0.0,5691,0,Camp Nelson,0,0,Fiber Optic,36.057458000000004,-118.591951,1,40.9,1,6,None,191,1,0,1,0,35,0,415.0,0.0,0.0,1383.6,0,0,93208
5602,1,0,0,0,6,1,0,DSL,1,0,1,1,Two year,1,Mailed check,80.25,493.4,0,50,10,22.95,2706,0,Coalinga,1,1,Fiber Optic,36.186867,-120.38779299999999,0,80.25,0,0,Offer E,18036,1,0,0,1,6,1,49.0,137.7,0.0,493.4,0,0,93210
5603,0,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),48.6,48.6,1,22,57,6.54,4207,1,Corcoran,0,0,DSL,36.04533,-119.532424,0,50.544,0,0,Offer E,23506,0,0,0,0,1,1,0.0,6.54,0.0,48.6,1,0,93212
5604,1,0,0,0,17,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.8,1207,0,26,52,35.88,5420,0,Delano,0,1,Fiber Optic,35.772244,-119.20968899999998,0,70.8,0,0,Offer D,37280,0,0,0,0,17,0,628.0,609.96,0.0,1207.0,1,0,93215
5605,1,0,1,1,10,1,0,DSL,0,0,1,0,Month-to-month,0,Mailed check,60.2,563.5,0,50,12,19.77,5318,0,Ducor,1,1,DSL,35.846067,-119.00407299999999,1,60.2,2,5,Offer D,823,0,0,1,0,10,0,0.0,197.7,0.0,563.5,0,1,93218
5606,1,0,0,1,15,1,0,DSL,0,0,0,0,One year,0,Credit card (automatic),55.2,864.55,0,62,11,1.63,3608,0,Earlimart,1,1,Fiber Optic,35.858053999999996,-119.305858,0,55.2,2,0,Offer D,9318,1,0,0,0,15,1,9.51,24.45,0.0,864.55,0,1,93219
5607,0,1,0,0,40,0,No phone service,DSL,1,1,1,1,Month-to-month,1,Electronic check,55.8,2109.35,1,72,7,0.0,4272,1,Exeter,0,0,Fiber Optic,36.301689,-119.01823300000001,0,58.032,0,0,None,13333,0,0,0,1,40,4,0.0,0.0,0.0,2109.35,0,1,93221
5608,0,0,1,1,13,1,0,DSL,1,0,0,0,One year,0,Bank transfer (automatic),54.15,701.05,0,51,12,19.63,4977,0,Frazier Park,0,0,DSL,34.907911,-119.23428100000001,1,54.15,1,5,Offer D,1526,1,0,1,0,13,3,84.0,255.19,0.0,701.05,0,0,93222
5609,1,0,1,0,29,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.15,2265.25,1,29,52,26.03,5189,1,Farmersville,0,1,Cable,36.29878,-119.20102800000001,1,83.35600000000002,0,1,Offer C,8644,0,0,1,0,29,9,1178.0,754.87,0.0,2265.25,1,0,93223
5610,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.5,220.6,1,30,94,47.51,5948,1,Fellows,0,0,Cable,35.215731,-119.57013,0,78.52,0,0,Offer E,626,0,2,0,0,3,4,207.0,142.53,0.0,220.6,0,0,93224
5611,0,1,1,0,58,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),100.4,5749.8,0,72,28,47.34,4005,0,Frazier Park,0,0,Cable,34.827662,-118.999073,1,100.4,0,8,Offer B,4498,1,0,1,1,58,0,0.0,2745.7200000000007,0.0,5749.8,0,1,93225
5612,0,0,0,0,45,1,0,DSL,1,1,0,0,One year,1,Credit card (automatic),62.55,2796.45,0,48,8,8.4,2935,0,Glennville,0,0,Cable,35.735694,-118.738483,0,62.55,0,0,Offer B,296,1,1,0,0,45,1,0.0,378.0,0.0,2796.45,0,1,93226
5613,0,0,1,1,72,1,1,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),70.45,5165.7,0,52,19,6.85,4463,0,Hanford,1,0,DSL,36.292229999999996,-119.622676,1,70.45,1,8,Offer A,53204,1,0,1,0,72,1,0.0,493.2,0.0,5165.7,0,1,93230
5614,1,0,1,1,68,1,1,Fiber optic,1,1,0,0,One year,1,Bank transfer (automatic),85.5,5696.6,0,27,85,29.67,4380,0,Huron,0,1,Fiber Optic,36.217864,-120.08011699999999,1,85.5,1,1,None,6918,0,0,1,0,68,0,4842.0,2017.56,0.0,5696.6,1,0,93234
5615,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.2,20.2,1,28,0,10.98,5394,1,Ivanhoe,0,1,NA,36.385818,-119.22424299999999,0,20.2,0,0,Offer E,4517,0,0,0,0,1,2,0.0,10.98,0.0,20.2,1,0,93235
5616,0,0,1,1,38,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,54.5,2076.05,0,30,30,46.27,5499,0,Kernville,0,0,Fiber Optic,35.852892,-118.397782,1,54.5,3,5,None,1873,0,0,1,0,38,2,0.0,1758.2600000000002,0.0,2076.05,0,1,93238
5617,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.75,44.2,0,35,0,27.67,3976,0,Kettleman City,0,1,NA,35.996922999999995,-120.000951,0,20.75,0,0,None,1809,0,0,0,0,2,0,0.0,55.34,0.0,44.2,0,0,93239
5618,1,0,0,0,11,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,215.25,0,43,0,47.88,5597,0,Lake Isabella,0,1,NA,35.607875,-118.46631799999999,0,20.35,0,0,Offer D,5564,0,2,0,0,11,1,0.0,526.6800000000002,0.0,215.25,0,0,93240
5619,0,1,1,0,20,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),91.0,1859.5,0,65,2,38.85,3748,0,Lamont,0,0,Cable,35.245034999999994,-118.905553,1,91.0,0,2,None,15364,0,0,1,1,20,0,0.0,777.0,0.0,1859.5,0,1,93241
5620,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),104.8,7470.1,0,58,15,40.49,4165,0,Laton,1,1,Fiber Optic,36.444232,-119.71828500000001,1,104.8,0,4,None,2900,0,0,1,1,72,0,0.0,2915.28,0.0,7470.1,0,1,93242
5621,0,0,1,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.75,229.5,1,39,14,35.18,3972,1,Lebec,0,0,Cable,34.845861,-118.88516299999999,1,77.74000000000002,0,1,Offer E,1247,0,2,1,0,3,8,32.0,105.54,0.0,229.5,0,0,93243
5622,1,0,0,0,23,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,104.05,2470.1,1,49,2,16.28,5963,1,Lemon Cove,1,1,Fiber Optic,36.462671,-118.99729099999999,0,108.212,0,0,Offer D,293,1,1,0,1,23,3,49.0,374.44000000000005,0.0,2470.1,0,0,93244
5623,1,0,0,0,40,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,51.1,2092.9,0,26,73,34.49,3355,0,Lemoore,0,1,DSL,36.303666,-119.825657,0,51.1,0,0,Offer B,30419,1,0,0,0,40,1,0.0,1379.6,0.0,2092.9,1,1,93245
5624,1,1,1,0,62,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Bank transfer (automatic),89.8,5629.55,0,65,3,27.49,4981,0,Lindsay,0,1,DSL,36.205465000000004,-119.085807,1,89.8,0,7,Offer B,15508,0,0,1,1,62,1,0.0,1704.38,0.0,5629.55,0,1,93247
5625,0,0,0,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.55,469.85,0,28,0,43.97,3169,0,Lost Hills,0,0,NA,35.637715,-119.893068,0,20.55,2,0,Offer D,2502,0,0,0,0,22,2,0.0,967.34,0.0,469.85,1,0,93249
5626,0,0,0,0,11,1,0,DSL,1,0,0,1,Month-to-month,0,Bank transfer (automatic),64.05,733.95,0,19,52,40.96,4171,0,Mc Farland,1,0,DSL,35.666886,-119.18671699999999,0,64.05,0,0,Offer D,10781,0,0,0,1,11,0,0.0,450.56,0.0,733.95,1,1,93250
5627,1,1,1,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.85,485.25,0,68,13,6.81,2259,0,Mc Kittrick,0,1,Fiber Optic,35.38381,-119.73088500000001,1,74.85,0,2,None,302,0,1,1,0,7,1,0.0,47.67,0.0,485.25,0,1,93251
5628,0,0,0,0,13,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Electronic check,96.65,1244.5,1,28,45,17.02,2110,1,Temecula,0,0,Cable,33.507255,-117.029473,0,100.516,0,0,Offer D,46171,0,0,0,0,13,0,560.0,221.26,0.0,1244.5,1,0,92592
5629,1,1,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,20.05,1,69,0,19.87,3491,1,New Cuyama,0,1,NA,34.956577,-119.750142,0,20.05,0,0,Offer E,798,0,0,0,0,1,4,0.0,19.87,0.0,20.05,0,0,93254
5630,0,0,0,0,39,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,103.45,3994.45,1,52,31,34.74,4811,1,Temecula,1,0,Cable,33.507255,-117.029473,0,107.588,0,0,Offer C,46171,0,0,0,1,39,1,1238.0,1354.86,0.0,3994.45,0,0,92592
5631,1,0,1,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,25.0,78.25,0,46,12,0.0,2730,0,Pixley,0,1,DSL,35.957019,-119.330928,1,25.0,0,1,Offer E,4198,0,0,1,0,3,1,9.0,0.0,0.0,78.25,0,0,93256
5632,1,0,0,0,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.3,1131.5,0,58,0,29.25,4335,0,Porterville,0,1,NA,36.008958,-118.891593,0,20.3,0,0,Offer B,65566,0,0,0,0,58,2,0.0,1696.5,0.0,1131.5,0,0,93257
5633,1,0,0,1,6,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,26.35,184.05,0,21,0,38.28,2189,0,Posey,0,1,NA,35.861928000000006,-118.636698,0,26.35,3,0,Offer E,266,0,0,0,0,6,0,0.0,229.68,0.0,184.05,1,0,93260
5634,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.9,19.9,1,33,0,7.49,4633,1,Richgrove,0,0,NA,35.809921,-119.12743700000001,1,19.9,1,1,None,2956,0,2,1,0,1,4,0.0,7.49,0.0,19.9,0,0,93261
5635,0,0,1,0,22,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,54.7,1178.75,0,60,16,39.83,5722,0,Sequoia National Park,1,0,DSL,36.527243,-118.59493799999998,1,54.7,0,1,Offer D,56,0,0,1,0,22,0,18.86,876.26,0.0,1178.75,0,1,93262
5636,1,0,1,0,14,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Electronic check,46.35,667.7,1,53,13,0.0,5360,1,Shafter,0,1,DSL,35.490705,-119.286833,1,48.20399999999999,0,1,Offer D,15177,0,1,1,1,14,4,0.0,0.0,0.0,667.7,0,1,93263
5637,1,0,1,1,64,1,1,Fiber optic,0,0,0,1,One year,0,Credit card (automatic),90.25,5629.15,0,57,30,45.35,4799,0,Springville,1,1,Fiber Optic,36.245926000000004,-118.69313799999999,1,90.25,2,9,Offer B,3546,0,0,1,1,64,0,1689.0,2902.4,0.0,5629.15,0,0,93265
5638,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.95,19.95,1,62,0,17.61,2051,1,Stratford,0,1,NA,36.175255,-119.813805,0,19.95,0,0,None,1729,0,2,0,0,1,2,0.0,17.61,0.0,19.95,0,0,93266
5639,1,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.65,109.3,0,33,0,32.34,3266,0,Strathmore,0,1,NA,36.141319,-119.129075,0,20.65,0,0,Offer E,5689,0,0,0,0,6,0,0.0,194.04,0.0,109.3,0,0,93267
5640,1,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,79.6,79.6,1,40,24,19.32,2199,1,Taft,0,1,DSL,35.184837,-119.402525,0,82.78399999999998,0,0,None,14937,0,0,0,1,1,5,0.0,19.32,0.0,79.6,0,0,93268
5641,1,0,0,1,39,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),25.45,958.45,0,45,0,46.57,5986,0,Terra Bella,0,1,NA,35.939068,-119.04366599999999,0,25.45,2,0,None,5868,0,0,0,0,39,0,0.0,1816.23,0.0,958.45,0,0,93270
5642,0,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.5,403.15,0,38,0,38.74,4700,0,Three Rivers,0,0,NA,36.413433000000005,-118.854708,0,19.5,0,0,None,2318,0,0,0,0,20,0,0.0,774.8000000000002,0.0,403.15,0,0,93271
5643,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.9,75.9,1,23,30,44.56,3389,1,Temecula,0,1,Fiber Optic,33.507255,-117.029473,0,78.936,0,0,None,46171,1,0,0,0,1,0,0.0,44.56,0.0,75.9,1,0,92592
5644,1,0,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,76.2,76.2,1,53,15,35.15,5973,1,Tulare,1,1,Fiber Optic,36.185471,-119.375243,1,79.248,0,1,None,56101,0,0,1,0,1,3,0.0,35.15,0.0,76.2,0,0,93274
5645,1,0,1,0,64,1,1,DSL,1,0,1,0,One year,1,Credit card (automatic),66.15,4392.5,0,40,2,37.46,4703,0,Tupman,0,1,Fiber Optic,35.316263,-119.40255900000001,1,66.15,0,3,Offer B,236,0,0,1,0,64,0,0.0,2397.44,0.0,4392.5,0,1,93276
5646,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.25,19.25,1,35,0,12.81,5437,1,Visalia,0,1,NA,36.303793,-119.375646,0,19.25,7,0,None,44741,0,2,0,0,1,4,0.0,12.81,0.0,19.25,0,0,93277
5647,0,0,1,0,46,1,0,DSL,0,1,1,1,Month-to-month,1,Credit card (automatic),69.1,3168,0,29,53,31.88,2333,0,Wasco,0,0,Fiber Optic,35.652242,-119.4464,1,69.1,0,7,Offer B,22760,0,0,1,1,46,0,0.0,1466.48,0.0,3168.0,1,1,93280
5648,0,1,1,1,28,0,No phone service,DSL,0,1,0,1,One year,1,Electronic check,39.1,1096.6,0,76,21,0.0,2305,0,Weldon,0,0,DSL,35.556470000000004,-118.244914,1,39.1,3,2,None,1935,0,0,1,1,28,0,230.0,0.0,0.0,1096.6,0,0,93283
5649,0,0,1,0,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,669.45,0,34,0,4.15,5759,0,Wofford Heights,0,0,NA,35.690535,-118.552784,1,20.05,0,5,None,2515,0,0,1,0,33,0,0.0,136.95000000000002,0.0,669.45,0,0,93285
5650,1,0,1,1,39,1,0,DSL,1,1,0,0,One year,0,Electronic check,59.8,2343.85,0,60,13,13.8,3093,0,Woodlake,1,1,Cable,36.464634999999994,-119.094348,1,59.8,2,5,None,8870,0,0,1,0,39,2,305.0,538.2,0.0,2343.85,0,0,93286
5651,0,0,1,0,42,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,84.3,3588.4,1,58,24,10.73,2514,1,Woody,1,0,DSL,35.710244,-118.881679,1,87.67200000000001,0,1,None,88,1,0,1,0,42,3,861.0,450.66,0.0,3588.4,0,0,93287
5652,0,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,48.6,48.6,0,51,11,7.99,3704,0,Visalia,0,0,Fiber Optic,36.391777000000005,-119.37284199999999,0,48.6,0,0,Offer E,36718,0,0,0,0,1,0,0.0,7.99,0.0,48.6,0,1,93291
5653,0,0,0,0,7,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.0,522.95,1,63,2,26.09,3735,1,Visalia,0,0,Fiber Optic,36.37559,-119.21168899999999,0,82.16,0,0,None,30395,0,1,0,0,7,2,10.0,182.63,0.0,522.95,0,0,93292
5654,1,1,1,0,70,1,0,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),105.35,7511.9,0,70,7,14.48,5866,0,Bakersfield,1,1,DSL,35.383937,-119.02042800000001,1,105.35,0,2,Offer A,12963,0,1,1,1,70,2,0.0,1013.6,0.0,7511.9,0,1,93301
5655,1,0,0,0,65,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.1,1725,0,22,0,20.43,5449,0,Bakersfield,0,1,NA,35.339796,-119.023552,0,25.1,0,0,Offer B,44588,0,0,0,0,65,0,0.0,1327.95,0.0,1725.0,1,0,93304
5656,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,49.75,49.75,0,47,14,41.79,2908,0,Bakersfield,0,1,Cable,35.391733,-118.984109,0,49.75,0,0,Offer E,35643,0,0,0,0,1,0,0.0,41.79,0.0,49.75,0,0,93305
5657,1,0,1,0,18,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.75,1691.9,0,42,16,34.17,4477,0,Bakersfield,0,1,Fiber Optic,35.449881,-118.84144199999999,1,94.75,0,1,None,53481,0,0,1,1,18,0,271.0,615.0600000000002,0.0,1691.9,0,0,93306
5658,1,0,1,0,24,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.0,2248.05,0,54,20,46.91,5886,0,Bakersfield,0,1,Fiber Optic,35.280113,-118.962329,1,93.0,0,7,None,59195,0,0,1,1,24,0,0.0,1125.84,0.0,2248.05,0,1,93307
5659,1,0,0,0,63,1,1,DSL,1,0,0,1,Two year,1,Bank transfer (automatic),71.9,4479.2,0,20,85,42.59,5816,0,Bakersfield,1,1,Cable,35.559616999999996,-118.92518500000001,0,71.9,0,0,Offer B,44915,1,0,0,1,63,1,3807.0,2683.17,0.0,4479.2,1,0,93308
5660,0,0,0,1,44,1,1,DSL,0,1,1,1,One year,1,Mailed check,77.55,3471.1,0,39,26,5.07,5044,0,Bakersfield,0,0,Fiber Optic,35.342890999999995,-119.064803,0,77.55,3,0,Offer B,58632,0,0,0,1,44,1,0.0,223.08,0.0,3471.1,0,1,93309
5661,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.85,63,0,26,0,6.88,5918,0,Bakersfield,0,1,NA,35.16207,-119.19448799999999,0,19.85,0,0,Offer E,20440,0,0,0,0,4,1,0.0,27.52,0.0,63.0,1,0,93311
5662,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.25,70.25,1,27,65,23.0,4133,1,Bakersfield,0,0,Fiber Optic,35.392599,-119.245341,0,73.06,0,0,Offer E,40836,0,4,0,0,1,3,0.0,23.0,0.0,70.25,1,0,93312
5663,0,0,1,1,37,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.25,3314.15,0,43,11,1.6,2969,0,Bakersfield,0,0,Fiber Optic,35.140938,-119.051348,1,95.25,2,0,None,25126,0,0,0,1,37,0,365.0,59.2,0.0,3314.15,0,0,93313
5664,0,1,0,0,10,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),84.6,865.55,1,70,33,16.85,3320,1,San Luis Obispo,1,0,Cable,35.233745,-120.626442,0,87.984,0,0,None,27047,0,0,0,1,10,6,286.0,168.5,0.0,865.55,0,0,93401
5665,1,0,0,0,34,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),25.05,852.7,0,59,28,0.0,3800,0,Los Osos,0,1,Fiber Optic,35.279984000000006,-120.824288,0,25.05,0,0,None,14859,0,0,0,0,34,2,239.0,0.0,0.0,852.7,0,0,93402
5666,1,0,1,0,35,0,No phone service,DSL,1,0,1,1,One year,0,Credit card (automatic),53.15,1930.9,0,53,30,0.0,5638,0,San Luis Obispo,1,1,DSL,35.236549,-120.72734399999999,1,53.15,0,5,None,31982,0,0,1,1,35,1,0.0,0.0,0.0,1930.9,0,1,93405
5667,0,0,1,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,20.15,91.4,0,35,0,45.84,2198,0,Arroyo Grande,0,0,NA,35.176235999999996,-120.48324299999999,1,20.15,0,5,None,24499,0,0,1,0,4,0,0.0,183.36,0.0,91.4,0,0,93420
5668,0,1,1,0,39,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.25,3949.15,0,73,21,20.15,3172,0,Atascadero,0,0,Cable,35.453912,-120.69461000000001,1,101.25,0,9,None,29539,1,0,1,1,39,0,829.0,785.8499999999998,0.0,3949.15,0,0,93422
5669,1,1,1,0,43,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),100.55,4304,0,77,8,37.09,4499,0,Avila Beach,1,1,Fiber Optic,35.186644,-120.728305,1,100.55,0,10,Offer B,812,0,2,1,1,43,2,344.0,1594.87,0.0,4304.0,0,0,93424
5670,0,0,1,1,17,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,24.1,409.9,1,31,0,18.26,4648,1,Bradley,0,0,NA,35.842889,-121.00486200000002,1,24.1,2,1,Offer D,1363,0,1,1,0,17,2,0.0,310.42,0.0,409.9,0,0,93426
5671,0,0,1,0,61,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.3,1554.9,0,52,0,40.37,4501,0,Buellton,0,0,NA,34.631362,-120.23821799999999,1,25.3,0,1,Offer B,4644,0,0,1,0,61,1,0.0,2462.57,0.0,1554.9,0,0,93427
5672,0,0,1,0,49,1,1,DSL,1,1,0,1,One year,0,Electronic check,71.8,3472.05,0,47,30,25.1,6193,0,Cambria,1,0,DSL,35.591387,-121.032256,1,71.8,0,9,Offer B,6526,0,0,1,1,49,1,0.0,1229.9,0.0,3472.05,0,1,93428
5673,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.7,117.8,0,49,0,23.04,5018,0,Casmalia,0,1,NA,34.866032000000004,-120.536546,0,19.7,0,0,None,210,0,0,0,0,4,0,0.0,92.16,0.0,117.8,0,0,93429
5674,0,0,1,1,64,0,No phone service,DSL,0,1,0,1,Two year,0,Electronic check,49.85,3210.35,0,28,59,0.0,5644,0,Cayucos,1,0,Cable,35.511833,-120.91871299999998,1,49.85,3,3,Offer B,3220,1,0,1,1,64,1,1894.0,0.0,0.0,3210.35,1,0,93430
5675,1,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.6,207.4,0,43,16,28.97,5487,0,Creston,0,1,Fiber Optic,35.480896,-120.469476,0,69.6,0,0,None,1203,0,0,0,0,3,0,33.0,86.91,0.0,207.4,0,0,93432
5676,1,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.75,19.75,0,31,0,30.38,3068,0,Grover Beach,0,1,NA,35.120833000000005,-120.61843,1,19.75,2,8,None,13106,0,0,1,0,1,0,0.0,30.38,0.0,19.75,0,0,93433
5677,1,0,1,0,40,1,0,Fiber optic,0,1,0,0,One year,0,Electronic check,80.8,3132.75,0,46,24,12.97,3387,0,Guadalupe,1,1,Fiber Optic,34.936,-120.594655,1,80.8,0,5,Offer B,5726,0,1,1,0,40,2,0.0,518.8000000000002,0.0,3132.75,0,1,93434
5678,0,0,0,1,1,1,0,DSL,1,1,0,0,Month-to-month,1,Electronic check,60.0,60,1,64,18,43.48,4531,1,Lompoc,0,0,Fiber Optic,34.601055,-120.38291699999999,0,62.40000000000001,2,0,Offer E,51737,1,1,0,0,1,2,0.0,43.48,0.0,60.0,0,0,93436
5679,1,0,0,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.55,649.65,1,47,2,24.76,4193,1,Lompoc,0,1,Cable,34.757477,-120.55050700000001,0,90.012,0,0,Offer E,6165,0,0,0,1,8,2,13.0,198.08,0.0,649.65,0,0,93437
5680,0,1,1,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.85,20.85,1,80,0,22.86,3817,1,Los Alamos,0,0,NA,34.758699,-120.27583899999999,1,20.85,0,1,Offer E,1328,0,0,1,0,1,2,0.0,22.86,0.0,20.85,0,0,93440
5681,0,1,1,0,34,1,0,DSL,0,0,1,0,One year,0,Bank transfer (automatic),64.2,2106.3,0,74,23,12.33,2225,0,Los Olivos,1,0,Cable,34.70434,-120.02609,1,64.2,0,2,None,1317,1,0,1,0,34,1,48.44,419.22,0.0,2106.3,0,1,93441
5682,0,0,1,0,1,0,No phone service,DSL,0,0,0,1,Month-to-month,0,Electronic check,35.0,35,0,33,14,0.0,4099,0,Morro Bay,0,0,Fiber Optic,35.369553,-120.76386399999998,1,35.0,0,9,None,10909,0,0,1,1,1,1,0.0,0.0,0.0,35.0,0,0,93442
5683,0,0,0,0,39,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,50.75,2011.4,1,35,4,0.0,4119,1,Nipomo,1,0,Cable,35.050345,-120.489599,0,52.78,0,0,Offer C,15405,0,0,0,1,39,6,80.0,0.0,0.0,2011.4,0,0,93444
5684,0,1,1,0,58,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),105.5,6205.5,1,73,21,16.94,5067,1,Oceano,0,0,Cable,35.059695,-120.60474099999999,1,109.72,0,1,None,7435,1,1,1,1,58,2,1303.0,982.52,0.0,6205.5,0,0,93445
5685,1,0,1,1,45,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Electronic check,19.2,903.7,0,21,0,17.23,3451,0,Paso Robles,0,1,NA,35.634221999999994,-120.72834099999999,1,19.2,1,6,Offer B,35586,0,0,1,0,45,1,0.0,775.35,0.0,903.7,1,0,93446
5686,1,1,0,0,6,1,0,Fiber optic,1,0,1,0,Month-to-month,1,Bank transfer (automatic),85.15,503.6,1,73,33,29.41,5831,1,Pismo Beach,0,1,DSL,35.165668,-120.65584199999999,0,88.55600000000003,0,0,Offer E,8564,0,0,0,0,6,4,166.0,176.46,0.0,503.6,0,0,93449
5687,1,0,0,0,43,1,0,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),90.65,3882.3,0,19,59,36.78,2496,0,San Ardo,1,1,DSL,35.996008,-120.85305,0,90.65,0,0,Offer B,670,1,0,0,0,43,1,2291.0,1581.54,0.0,3882.3,1,0,93450
5688,1,0,1,1,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.0,879.8,0,24,0,16.02,5743,0,San Miguel,0,1,NA,35.886767,-120.60866100000001,1,20.0,1,5,None,2666,0,0,1,0,41,0,0.0,656.8199999999998,0.0,879.8,1,0,93451
5689,1,0,0,0,5,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.65,383.65,0,58,16,32.81,3319,0,San Simeon,0,1,DSL,35.746484,-121.223355,0,74.65,0,0,None,471,0,0,0,0,5,1,6.14,164.05,0.0,383.65,0,1,93452
5690,1,0,0,0,72,0,No phone service,DSL,1,0,1,1,Two year,1,Credit card (automatic),61.2,4390.25,0,43,6,0.0,4085,0,Santa Margarita,1,1,Cable,35.303926000000004,-120.25656699999999,0,61.2,0,0,None,2687,1,0,0,1,72,0,0.0,0.0,0.0,4390.25,0,1,93453
5691,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.95,68.2,0,47,0,6.86,2195,0,Santa Maria,0,1,NA,34.943523,-120.256729,0,19.95,0,0,None,30540,0,0,0,0,4,1,0.0,27.44,0.0,68.2,0,0,93454
5692,1,0,1,1,9,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,54.8,452.8,0,43,24,44.46,2848,0,Santa Maria,0,1,DSL,34.818227,-120.418784,1,54.8,2,2,None,37364,1,1,1,0,9,1,0.0,400.14,0.0,452.8,0,1,93455
5693,1,1,1,0,72,1,1,DSL,0,0,1,1,Two year,1,Credit card (automatic),73.45,5329,0,79,3,11.26,5540,0,Santa Maria,1,1,DSL,34.959340000000005,-120.490081,1,73.45,0,7,Offer A,43684,0,0,1,1,72,2,15.99,810.72,0.0,5329.0,0,1,93458
5694,0,0,1,0,33,1,0,DSL,0,0,0,0,One year,1,Mailed check,51.45,1758.9,0,42,9,48.09,4935,0,Santa Ynez,0,0,Cable,34.630356,-120.032564,1,51.45,0,7,None,5710,1,0,1,0,33,0,158.0,1586.97,0.0,1758.9,0,0,93460
5695,0,0,1,0,72,1,1,Fiber optic,1,0,0,0,Two year,0,Bank transfer (automatic),80.45,5737.6,0,59,27,6.23,4202,0,Shandon,0,0,Fiber Optic,35.634488,-120.29353400000001,1,80.45,0,4,None,1255,0,0,1,0,72,1,1549.0,448.56000000000006,0.0,5737.6,0,0,93461
5696,1,0,1,0,22,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,54.2,1152.7,1,48,23,27.24,5102,1,Solvang,0,1,DSL,34.624399,-120.137875,1,56.368,0,1,Offer D,7958,1,0,1,0,22,3,265.0,599.28,0.0,1152.7,0,0,93463
5697,0,0,1,0,70,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,109.5,7674.55,1,21,65,41.88,4191,1,Templeton,1,0,DSL,35.536115,-120.739231,1,113.88,0,1,Offer A,7918,1,0,1,1,70,2,4988.0,2931.600000000001,0.0,7674.55,1,0,93465
5698,1,0,1,1,21,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,104.4,2157.95,1,45,3,42.65,3796,1,Mojave,1,1,DSL,35.097322999999996,-118.17128799999999,1,108.576,0,1,Offer D,4882,0,0,1,1,21,5,6.47,895.65,0.0,2157.95,0,1,93501
5699,1,0,0,0,15,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,85.3,1219.85,0,41,18,27.3,5559,0,California City,1,1,Fiber Optic,35.151491,-117.92759699999999,0,85.3,0,0,None,8316,0,0,0,0,15,0,0.0,409.5,0.0,1219.85,0,1,93505
5700,1,1,1,0,29,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,79.3,2414.55,0,69,2,10.55,3172,0,Acton,0,1,Fiber Optic,34.501452,-118.207862,1,79.3,0,0,None,7831,1,0,0,0,29,0,0.0,305.9500000000001,0.0,2414.55,0,1,93510
5701,0,0,1,1,15,1,0,DSL,0,1,1,1,Month-to-month,0,Bank transfer (automatic),76.5,1155.6,0,63,18,39.77,3851,0,Benton,1,0,Cable,37.653946999999995,-118.231443,1,76.5,1,5,None,340,1,0,1,1,15,0,20.8,596.5500000000002,0.0,1155.6,0,1,93512
5702,1,1,1,1,71,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),105.1,7548.1,1,79,9,44.66,5725,1,Big Pine,0,1,DSL,37.245505,-118.06294299999999,1,109.304,0,1,None,1826,0,1,1,1,71,3,679.0,3170.86,0.0,7548.1,0,0,93513
5703,1,1,0,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.4,1809.35,0,80,0,26.01,6141,0,Bishop,0,1,NA,37.045840000000005,-118.397236,0,25.4,0,0,Offer A,13309,0,0,0,0,72,1,0.0,1872.72,0.0,1809.35,0,0,93514
5704,0,0,1,0,19,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.85,1564.4,0,34,16,7.84,5072,0,Boron,0,0,Fiber Optic,34.957029999999996,-117.73045,1,86.85,0,8,None,2241,0,0,1,0,19,1,250.0,148.96,0.0,1564.4,0,0,93516
5705,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,19.65,0,40,0,16.91,3192,0,Bridgeport,0,1,NA,38.184583,-119.28655800000001,0,19.65,0,0,None,826,0,1,0,0,1,1,0.0,16.91,0.0,19.65,0,0,93517
5706,0,0,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,75.7,75.7,1,39,23,9.05,4884,1,Caliente,0,0,Fiber Optic,35.358953,-118.527064,0,78.72800000000002,0,0,Offer E,1022,0,0,0,0,1,4,0.0,9.05,0.0,75.7,0,0,93518
5707,0,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.55,84.4,0,26,71,41.9,4372,0,Darwin,0,0,Fiber Optic,36.319181,-117.593053,0,45.55,0,0,Offer E,64,0,0,0,0,2,0,0.0,83.8,0.0,84.4,1,1,93522
5708,0,1,1,1,11,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),78.1,864.85,0,77,13,17.66,2333,0,Edwards,1,0,Cable,34.966777,-117.961179,1,78.1,2,8,None,7685,0,0,1,0,11,0,0.0,194.26,0.0,864.85,0,1,93523
5709,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.3,228.75,0,58,0,41.78,2868,0,Independence,0,0,NA,36.869584,-118.189241,0,19.3,0,0,None,734,0,0,0,0,12,0,0.0,501.36,0.0,228.75,0,0,93526
5710,0,0,1,0,70,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,110.5,7752.05,0,41,23,28.54,5979,0,Temecula,1,0,DSL,33.507255,-117.029473,1,110.5,0,4,None,46171,1,0,1,1,70,0,1783.0,1997.8,0.0,7752.05,0,0,92592
5711,0,1,1,0,20,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,90.8,1951,1,79,19,4.77,2312,1,Johannesburg,1,0,Cable,35.363339,-117.63764099999999,1,94.432,0,1,None,207,0,2,1,0,20,1,0.0,95.4,0.0,1951.0,0,1,93528
5712,0,0,0,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),20.3,470.6,0,38,0,16.26,3630,0,June Lake,0,0,NA,37.730269,-119.05581299999999,0,20.3,0,0,None,618,0,0,0,0,23,0,0.0,373.98,0.0,470.6,0,0,93529
5713,1,1,0,0,49,1,1,DSL,1,1,0,1,Two year,0,Credit card (automatic),81.35,4060.9,0,67,10,43.19,4537,0,Keeler,1,1,Fiber Optic,36.560497999999995,-117.962461,0,81.35,0,0,Offer B,71,1,0,0,1,49,1,406.0,2116.31,0.0,4060.9,0,0,93530
5714,0,0,1,1,4,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,97.95,384.5,1,21,56,9.98,2570,1,Keene,0,0,Cable,35.214982,-118.59048999999999,1,101.868,0,4,Offer E,1436,0,0,1,1,4,4,215.0,39.92,0.0,384.5,1,0,93531
5715,1,0,0,0,32,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Credit card (automatic),108.15,3432.9,1,22,80,27.69,2541,1,Lake Hughes,0,1,DSL,34.659579,-118.58421200000001,0,112.476,0,0,Offer C,2771,1,0,0,1,32,3,2746.0,886.08,0.0,3432.9,1,0,93532
5716,1,0,0,1,2,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.3,108.65,0,22,59,43.93,4594,0,Lancaster,0,1,DSL,34.727529,-118.153098,0,55.3,1,0,Offer E,35109,0,0,0,1,2,0,64.0,87.86,0.0,108.65,1,0,93534
5717,1,1,1,0,69,0,No phone service,DSL,1,1,1,1,Two year,0,Credit card (automatic),56.55,3952.65,0,79,12,0.0,4162,0,Lancaster,0,1,DSL,34.712708,-117.889656,1,56.55,0,10,Offer A,57794,0,0,1,1,69,0,474.0,0.0,0.0,3952.65,0,0,93535
5718,1,0,0,0,6,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),80.5,463.05,1,45,29,6.4,2181,1,Lancaster,0,1,Fiber Optic,34.741406,-118.38111,0,83.72,0,0,None,49309,0,0,0,0,6,1,0.0,38.40000000000001,0.0,463.05,0,1,93536
5719,0,0,1,1,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.7,494.05,0,43,0,46.3,3594,0,Lee Vining,0,0,NA,37.890145000000004,-119.184087,1,19.7,3,5,None,504,0,0,1,0,24,2,0.0,1111.1999999999996,0.0,494.05,0,0,93541
5720,0,0,0,0,32,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),104.05,3416.85,0,44,28,14.21,2335,0,Littlerock,1,0,Fiber Optic,34.505272999999995,-117.955054,0,104.05,0,0,None,11198,0,0,0,1,32,0,957.0,454.72,0.0,3416.85,0,0,93543
5721,0,0,0,0,27,1,0,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),52.85,1498.65,0,44,29,10.55,2842,0,Llano,0,0,Fiber Optic,34.500091,-117.76586200000001,0,52.85,0,0,None,1220,0,0,0,0,27,2,0.0,284.85,0.0,1498.65,0,1,93544
5722,0,1,1,0,27,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Bank transfer (automatic),104.3,2867.75,1,73,30,10.19,3444,1,Fallbrook,0,0,Fiber Optic,33.362575,-117.299644,1,108.47200000000001,0,5,Offer C,42239,1,0,1,0,27,2,860.0,275.13,0.0,2867.75,0,0,92028
5723,1,0,0,0,58,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),80.65,4807.35,0,52,8,44.67,6043,0,Mammoth Lakes,0,1,DSL,37.550074,-118.837167,0,80.65,0,0,None,8217,1,0,0,0,58,0,385.0,2590.86,0.0,4807.35,0,0,93546
5724,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,71.35,71.35,1,23,56,35.28,5730,1,Olancha,0,1,Cable,36.296851000000004,-117.86546899999999,0,74.204,0,0,None,318,0,0,0,1,1,5,0.0,35.28,0.0,71.35,1,0,93549
5725,0,0,1,1,18,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.65,471.35,0,22,0,43.69,5231,0,Palmdale,0,0,NA,34.536232,-118.082935,1,24.65,3,9,None,67232,0,0,1,0,18,2,0.0,786.42,0.0,471.35,1,0,93550
5726,0,0,1,1,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),21.3,1041.8,0,47,0,3.95,2861,0,Palmdale,0,0,NA,34.613476,-118.256358,1,21.3,3,5,None,34045,0,0,1,0,47,0,0.0,185.65,0.0,1041.8,0,0,93551
5727,0,0,1,1,70,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,110.2,7689.8,0,26,85,5.51,4098,0,Palmdale,1,0,DSL,34.557711,-118.02944099999999,1,110.2,3,4,None,25370,1,0,1,1,70,0,0.0,385.7,0.0,7689.8,1,1,93552
5728,0,0,0,0,13,1,1,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,89.4,1132.35,1,42,16,8.59,2226,1,Pearblossom,1,0,Cable,34.445239,-117.89486799999999,0,92.976,0,0,Offer D,1613,1,1,0,0,13,2,0.0,111.67,0.0,1132.35,0,1,93553
5729,0,0,1,1,36,1,0,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),51.05,1815,0,32,19,19.73,2161,0,Randsburg,0,0,DSL,35.405722,-117.773354,1,51.05,2,3,None,117,0,0,1,0,36,0,345.0,710.28,0.0,1815.0,0,0,93554
5730,1,0,0,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.8,1311.3,0,31,0,4.72,4260,0,Temecula,0,1,NA,33.507255,-117.029473,0,19.8,0,0,None,46171,0,0,0,0,67,0,0.0,316.24,0.0,1311.3,0,0,92592
5731,0,0,0,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.9,199.45,0,56,0,23.84,5811,0,Rosamond,0,0,NA,34.903052,-118.41125100000001,0,19.9,0,0,None,14931,0,0,0,0,10,1,0.0,238.4,0.0,199.45,0,0,93560
5732,1,1,0,0,19,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,87.3,1637.3,0,66,16,29.8,4447,0,Tehachapi,0,1,DSL,35.073777,-118.65211200000002,0,87.3,0,0,None,25805,0,0,0,1,19,1,0.0,566.2,0.0,1637.3,0,1,93561
5733,0,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.85,1326.35,0,43,0,16.84,6342,0,Temecula,0,0,NA,33.507255,-117.029473,1,19.85,2,2,None,46171,0,0,1,0,71,0,0.0,1195.64,0.0,1326.35,0,0,92592
5734,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Mailed check,89.4,6376.55,0,45,19,2.75,6044,0,Valyermo,1,1,DSL,34.39583,-117.734568,1,89.4,2,7,None,413,1,0,1,1,72,1,1212.0,198.0,0.0,6376.55,0,0,93563
5735,0,0,1,1,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.0,935.9,0,19,0,9.77,2608,0,Palmdale,0,0,NA,34.598221,-117.79593,1,20.0,3,2,None,6787,0,0,1,0,48,0,0.0,468.96,0.0,935.9,1,0,93591
5736,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,20.05,0,56,0,13.51,2067,0,Ahwahnee,0,1,NA,37.375816,-119.739935,0,20.05,0,0,None,1968,0,0,0,0,1,2,0.0,13.51,0.0,20.05,0,0,93601
5737,1,0,1,1,18,1,0,DSL,1,0,1,1,Month-to-month,0,Electronic check,83.25,1611.15,0,29,59,10.29,2065,0,Auberry,1,1,DSL,36.991762,-119.242874,1,83.25,1,3,None,3464,1,0,1,1,18,1,0.0,185.22,0.0,1611.15,1,1,93602
5738,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.6,20.6,1,56,0,47.26,3618,1,Badger,0,1,NA,36.64545,-118.924982,0,20.6,0,0,Offer E,273,0,0,0,0,1,1,0.0,47.26,0.0,20.6,0,0,93603
5739,1,1,1,0,67,1,1,Fiber optic,0,1,1,1,Two year,0,Bank transfer (automatic),102.9,6989.7,0,72,17,48.68,5869,0,Bass Lake,0,1,Fiber Optic,37.458366999999996,-119.34501100000001,1,102.9,0,9,Offer A,613,1,0,1,1,67,3,1188.0,3261.56,0.0,6989.7,0,0,93604
5740,1,0,1,1,69,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,39.1,2779.5,0,52,11,0.0,5987,0,Big Creek,1,1,Fiber Optic,37.17277,-119.2997,1,39.1,1,3,None,273,1,1,1,0,69,2,0.0,0.0,0.0,2779.5,0,1,93605
5741,1,0,0,0,19,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.95,1931.75,1,54,20,2.19,3670,1,Biola,0,1,Cable,36.798882,-120.01951100000001,0,103.948,0,0,Offer D,807,0,2,0,1,19,2,386.0,41.61,0.0,1931.75,0,0,93606
5742,1,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Mailed check,114.5,8331.95,0,75,19,5.6,6051,0,Cantua Creek,1,1,Fiber Optic,36.488056,-120.40769099999999,1,114.5,0,4,Offer A,1766,1,1,1,1,72,2,1583.0,403.2,0.0,8331.95,0,0,93608
5743,0,1,0,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.2,735.9,0,65,0,4.09,4947,0,Caruthers,0,0,NA,36.5276,-119.865999,0,20.2,0,0,None,5446,0,0,0,0,38,0,0.0,155.42,0.0,735.9,0,0,93609
5744,1,1,1,0,40,1,0,DSL,0,0,0,1,One year,0,Electronic check,55.8,2283.3,0,71,18,28.56,3587,0,Chowchilla,0,1,Cable,37.100947999999995,-120.27013600000001,1,55.8,0,8,None,19391,0,0,1,1,40,1,0.0,1142.4,0.0,2283.3,0,1,93610
5745,0,0,1,1,61,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.2,1445.2,0,56,0,34.84,6201,0,Clovis,0,0,NA,36.917652000000004,-119.59375700000001,1,24.2,1,7,None,46858,0,0,1,0,61,0,0.0,2125.24,0.0,1445.2,0,0,93611
5746,0,0,0,0,10,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),81.0,818.05,1,46,21,49.5,2946,1,Clovis,0,0,DSL,36.814539,-119.711868,0,84.24000000000002,0,0,Offer D,33856,0,0,0,0,10,1,172.0,495.0,0.0,818.05,0,0,93612
5747,1,0,1,0,32,1,1,DSL,1,0,1,0,One year,1,Credit card (automatic),72.8,2333.05,0,26,46,15.41,3278,0,Coarsegold,0,1,Cable,37.212191,-119.749323,1,72.8,0,10,None,9395,1,1,1,0,32,2,0.0,493.12,0.0,2333.05,1,1,93614
5748,0,0,0,0,21,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),99.85,1992.55,0,24,48,24.86,2113,0,Cutler,0,0,DSL,36.497895,-119.28548400000001,0,99.85,0,0,None,5519,0,0,0,1,21,1,956.0,522.06,0.0,1992.55,1,0,93615
5749,0,1,0,0,59,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,99.5,5890,0,70,9,24.27,5513,0,Del Rey,1,0,Fiber Optic,36.657462,-119.595293,0,99.5,0,0,None,1965,0,1,0,1,59,1,530.0,1431.93,0.0,5890.0,0,0,93616
5750,0,1,1,0,13,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.15,916.75,1,77,21,37.86,5101,1,Dinuba,0,0,Cable,36.523619000000004,-119.38686799999999,1,72.956,0,2,None,24206,0,1,1,0,13,3,0.0,492.18,0.0,916.75,0,1,93618
5751,0,0,0,0,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.25,1029.8,0,50,0,8.85,5134,0,Dos Palos,0,0,NA,37.045728000000004,-120.63068200000001,0,20.25,0,0,None,9388,0,0,0,0,47,1,0.0,415.95,0.0,1029.8,0,0,93620
5752,1,0,1,1,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),26.0,1796.55,0,63,0,11.6,4933,0,Dunlap,0,1,NA,36.789213000000004,-119.14033799999999,1,26.0,2,5,None,506,0,0,1,0,69,0,0.0,800.4,0.0,1796.55,0,0,93621
5753,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.9,33.7,0,56,0,3.82,5824,0,Firebaugh,0,1,NA,36.785618,-120.625382,0,19.9,0,0,Offer E,9491,0,0,0,0,2,2,0.0,7.64,0.0,33.7,0,0,93622
5754,0,0,1,1,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.05,454.05,0,35,0,46.45,4312,0,Fish Camp,0,0,NA,37.483534999999996,-119.679414,1,19.05,1,0,Offer D,77,0,0,0,0,22,1,0.0,1021.9,0.0,454.05,0,0,93623
5755,1,1,1,0,15,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Electronic check,96.5,1392.25,0,79,26,22.83,2394,0,Five Points,1,1,Fiber Optic,36.397745,-120.11991100000002,1,96.5,0,9,None,1852,0,0,1,0,15,2,362.0,342.45,0.0,1392.25,0,0,93624
5756,0,0,0,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.85,1049.6,0,62,0,18.81,6338,0,Fowler,0,0,NA,36.625792,-119.67248300000001,0,19.85,0,0,None,5635,0,0,0,0,53,0,0.0,996.93,0.0,1049.6,0,0,93625
5757,0,1,1,0,28,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,25.7,734.6,0,79,0,25.57,3136,0,Friant,0,0,NA,37.027663000000004,-119.69056,1,25.7,0,8,None,1125,0,0,1,0,28,1,0.0,715.96,0.0,734.6,0,0,93626
5758,1,0,0,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.3,475.1,0,42,0,10.36,4510,0,Helm,0,1,NA,36.520537,-120.118055,0,20.3,0,0,Offer D,152,0,0,0,0,22,0,0.0,227.92,0.0,475.1,0,0,93627
5759,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.15,70.15,1,53,10,42.09,5773,1,Hume,0,0,Fiber Optic,36.807595,-118.901544,0,72.956,0,0,Offer E,93,0,1,0,0,1,2,0.0,42.09,0.0,70.15,0,1,93628
5760,1,1,1,0,16,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,91.55,1540.05,0,66,20,15.44,4045,0,Kerman,1,1,DSL,36.727418,-120.123526,1,91.55,0,1,None,14062,1,1,1,1,16,1,308.0,247.04,0.0,1540.05,0,0,93630
5761,0,0,1,1,48,0,No phone service,DSL,1,1,0,0,Two year,0,Mailed check,39.4,1978.65,0,29,52,0.0,5701,0,Kingsburg,0,0,DSL,36.478239,-119.52136999999999,1,39.4,3,5,None,14088,1,0,1,0,48,0,102.89,0.0,0.0,1978.65,1,1,93631
5762,1,1,1,0,30,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Bank transfer (automatic),105.7,3181.8,0,75,22,33.48,2455,0,Lakeshore,1,1,Fiber Optic,37.290606,-119.216328,1,105.7,0,6,None,52,1,2,1,0,30,2,0.0,1004.4,0.0,3181.8,0,1,93634
5763,0,0,0,0,3,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.25,229.7,0,33,10,25.4,2156,0,Los Banos,0,0,DSL,36.995162,-120.955099,0,70.25,0,0,Offer E,29124,0,2,0,0,3,1,23.0,76.19999999999997,0.0,229.7,0,0,93635
5764,1,1,0,0,57,1,1,Fiber optic,1,0,0,1,Two year,0,Electronic check,93.75,5625.55,0,77,11,2.21,4276,0,Madera,0,1,Fiber Optic,36.902954,-120.194274,0,93.75,0,0,None,28434,1,0,0,1,57,0,0.0,125.97,0.0,5625.55,0,1,93637
5765,0,1,1,0,68,1,1,Fiber optic,1,1,0,1,One year,1,Credit card (automatic),96.55,6581.9,1,68,21,1.98,5957,1,Madera,0,0,Cable,37.004068,-119.930027,1,100.412,0,5,None,49247,0,1,1,0,68,1,0.0,134.64,0.0,6581.9,0,1,93638
5766,0,0,1,0,23,1,0,DSL,0,0,1,0,One year,0,Bank transfer (automatic),60.0,1347.15,0,55,18,1.39,3835,0,Escondido,0,0,Fiber Optic,33.141265000000004,-116.967221,1,60.0,0,5,Offer D,48690,1,0,1,0,23,3,0.0,31.97,0.0,1347.15,0,1,92027
5767,0,0,1,0,65,1,0,DSL,0,0,1,0,Two year,1,Credit card (automatic),59.8,3808.2,0,46,14,10.23,6034,0,Miramonte,0,0,Fiber Optic,36.696759,-119.024051,1,59.8,0,7,None,571,1,0,1,0,65,0,533.0,664.95,0.0,3808.2,0,0,93641
5768,1,0,1,0,44,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),90.65,3974.15,0,30,53,23.75,3786,0,North Fork,0,1,Fiber Optic,37.244307,-119.470256,1,90.65,0,7,None,3376,0,0,1,1,44,0,0.0,1045.0,0.0,3974.15,0,1,93643
5769,0,0,1,1,71,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),109.0,7661.8,0,22,69,1.84,4204,0,Oakhurst,1,0,Fiber Optic,37.648647,-119.231447,1,109.0,1,2,None,8521,0,0,1,1,71,4,0.0,130.64,0.0,7661.8,1,1,93644
5770,0,0,1,0,37,1,1,DSL,1,0,0,0,One year,0,Credit card (automatic),68.1,2479.25,0,64,11,30.36,2873,0,O Neals,1,0,Fiber Optic,37.140104,-119.65709199999999,1,68.1,0,1,None,173,1,0,1,0,37,0,0.0,1123.32,0.0,2479.25,0,1,93645
5771,0,0,0,0,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,266.6,0,53,0,23.2,4497,0,Orange Cove,0,0,NA,36.633497999999996,-119.298895,0,20.4,0,0,Offer D,8449,0,0,0,0,12,0,0.0,278.4,0.0,266.6,0,0,93646
5772,1,0,1,1,69,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),81.95,5601.4,0,20,48,49.16,6182,0,Orosi,1,1,Cable,36.600184999999996,-119.175655,1,81.95,2,1,Offer A,9780,1,0,1,1,69,0,2689.0,3392.04,0.0,5601.4,1,0,93647
5773,0,0,0,0,35,1,0,DSL,1,1,0,0,Month-to-month,0,Electronic check,60.55,1982.6,0,57,20,44.81,3463,0,Parlier,1,0,Fiber Optic,36.622237,-119.521126,0,60.55,0,0,None,12587,0,0,0,0,35,2,0.0,1568.35,0.0,1982.6,0,1,93648
5774,1,0,0,0,5,1,0,DSL,0,1,0,1,Month-to-month,1,Bank transfer (automatic),65.6,339.9,0,22,59,8.6,5636,0,Fresno,0,1,Fiber Optic,36.841654999999996,-119.79711299999998,0,65.6,0,0,None,3258,1,1,0,1,5,1,0.0,43.0,0.0,339.9,1,1,93650
5775,1,0,1,1,58,1,1,Fiber optic,0,0,1,0,Two year,0,Bank transfer (automatic),82.5,4828.05,0,40,24,29.93,4348,0,Prather,0,1,DSL,37.007238,-119.505661,1,82.5,2,1,None,1314,0,0,1,0,58,1,1159.0,1735.94,0.0,4828.05,0,0,93651
5776,1,0,1,0,72,1,1,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),82.3,5980.55,0,56,30,29.29,5219,0,Raisin City,1,1,Cable,36.594542,-119.905245,1,82.3,0,1,Offer A,265,1,0,1,1,72,0,0.0,2108.88,0.0,5980.55,0,1,93652
5777,1,0,1,0,72,1,1,DSL,1,1,0,0,Two year,0,Mailed check,68.15,4808.7,0,56,17,17.31,4613,0,Raymond,1,1,DSL,37.252057,-119.95783,1,68.15,0,1,Offer A,972,1,0,1,0,72,0,817.0,1246.32,0.0,4808.7,0,0,93653
5778,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.3,20.3,0,48,0,4.09,2507,0,Reedley,0,0,NA,36.636638,-119.421842,0,20.3,0,0,None,25923,0,0,0,0,1,1,0.0,4.09,0.0,20.3,0,0,93654
5779,0,0,0,0,39,1,0,Fiber optic,1,0,1,0,One year,1,Electronic check,95.55,3692.85,1,29,78,4.48,2767,1,Riverdale,1,0,Cable,36.452211,-119.94575,0,99.37200000000001,0,0,Offer C,5729,1,0,0,1,39,0,288.04,174.72000000000003,0.0,3692.85,1,1,93656
5780,1,0,1,1,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.2,1068.15,0,38,0,20.44,6050,0,Sanger,0,1,NA,36.819628,-119.44041399999999,1,20.2,3,1,None,28991,0,0,1,0,53,0,0.0,1083.3200000000004,0.0,1068.15,0,0,93657
5781,0,0,0,0,27,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.2,2383.6,0,31,2,39.62,4384,0,San Joaquin,1,0,DSL,36.600193,-120.153393,0,89.2,0,0,Offer C,4318,1,0,0,1,27,1,0.0,1069.74,0.0,2383.6,0,1,93660
5782,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.65,69.65,1,70,6,31.13,4741,1,Selma,0,0,Cable,36.545322,-119.64228100000001,0,72.436,0,0,None,26213,0,0,0,0,1,0,0.0,31.13,0.0,69.65,0,0,93662
5783,0,1,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.3,89.3,1,68,33,30.23,3067,1,Shaver Lake,0,0,Cable,37.223,-119.001021,0,92.87200000000001,0,0,Offer E,642,0,3,0,0,1,1,0.0,30.23,0.0,89.3,0,0,93664
5784,0,0,1,0,18,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,74.8,1438.05,0,25,41,43.29,4809,0,South Dos Palos,0,0,Fiber Optic,36.959731,-120.65351899999999,1,74.8,0,1,Offer D,343,0,0,1,0,18,2,590.0,779.22,0.0,1438.05,1,0,93665
5785,1,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.2,917.45,0,54,0,45.92,3136,0,Sultana,0,1,NA,36.545353000000006,-119.33853500000001,1,20.2,1,1,None,306,0,0,1,0,46,0,0.0,2112.32,0.0,917.45,0,0,93666
5786,0,0,1,0,72,1,1,DSL,1,0,1,1,Two year,1,Credit card (automatic),84.4,6096.45,0,38,28,5.25,5046,0,Tollhouse,1,0,Fiber Optic,36.993666,-119.34826699999999,1,84.4,0,1,Offer A,2633,1,0,1,1,72,1,0.0,378.0,0.0,6096.45,0,1,93667
5787,0,0,0,0,36,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,87.55,3078.1,1,42,26,27.72,2558,1,Tranquillity,1,0,Cable,36.635661,-120.28864399999999,0,91.052,0,0,None,1130,1,1,0,1,36,4,800.0,997.92,0.0,3078.1,0,0,93668
5788,0,0,1,0,4,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,25.15,99.95,0,55,29,0.0,3891,0,Wishon,0,0,Fiber Optic,37.287758000000004,-119.548156,1,25.15,0,1,None,327,0,0,1,0,4,4,29.0,0.0,0.0,99.95,0,0,93669
5789,0,0,0,0,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.8,475.2,0,42,0,13.93,3875,0,Traver,0,0,NA,36.456091,-119.486225,0,19.8,0,0,Offer C,646,0,0,0,0,25,1,0.0,348.25,0.0,475.2,0,0,93673
5790,0,0,1,1,40,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,50.85,2036.55,0,27,52,0.0,2819,0,Squaw Valley,0,0,Fiber Optic,36.719141,-119.20267700000001,1,50.85,3,0,None,3146,0,1,0,1,40,1,1059.0,0.0,0.0,2036.55,1,0,93675
5791,1,0,1,0,63,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,102.4,6444.05,0,47,15,17.75,5096,0,Fresno,1,1,Fiber Optic,36.749403,-119.78757399999999,1,102.4,0,1,None,13858,0,0,1,1,63,1,967.0,1118.25,0.0,6444.05,0,0,93701
5792,0,1,0,0,15,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Mailed check,96.3,1426.75,1,76,9,19.11,2933,1,Fresno,1,0,Fiber Optic,36.739385,-119.753649,0,100.152,0,0,None,47999,1,0,0,0,15,6,128.0,286.65,0.0,1426.75,0,0,93702
5793,1,0,0,0,14,1,1,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),55.5,767.55,0,54,21,18.48,3520,0,Fresno,0,1,Fiber Optic,36.768774,-119.76263300000001,0,55.5,0,0,Offer D,31180,0,0,0,0,14,1,0.0,258.72,0.0,767.55,0,1,93703
5794,1,1,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),109.75,7932.5,0,66,14,18.74,4265,0,Fresno,1,1,Fiber Optic,36.799648,-119.801247,1,109.75,0,1,Offer A,26580,1,0,1,1,72,1,0.0,1349.28,0.0,7932.5,0,1,93704
5795,1,0,0,0,39,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,106.4,4040.65,0,55,30,17.17,4111,0,Fresno,0,1,DSL,36.787240000000004,-119.82781299999999,0,106.4,0,0,Offer C,35451,0,0,0,1,39,0,1212.0,669.6300000000001,0.0,4040.65,0,0,93705
5796,0,0,1,1,47,0,No phone service,DSL,1,1,1,1,Two year,1,Credit card (automatic),60.0,2768.65,0,37,25,0.0,3248,0,Fresno,1,0,Fiber Optic,36.654614,-119.903674,1,60.0,2,1,None,35790,0,0,1,1,47,0,69.22,0.0,0.0,2768.65,0,1,93706
5797,1,0,1,0,19,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),88.8,1672.35,0,42,20,34.05,4600,0,Fresno,0,1,DSL,36.822715,-119.761826,1,88.8,0,1,Offer D,29337,1,0,1,0,19,2,334.0,646.9499999999998,0.0,1672.35,0,0,93710
5798,0,0,0,0,5,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.2,474.8,1,26,51,34.49,4109,1,San Dimas,0,0,Fiber Optic,34.102119,-117.815532,0,88.60799999999999,0,0,Offer E,33878,0,0,0,1,5,6,242.0,172.45000000000005,0.0,474.8,1,0,91773
5799,0,0,0,0,13,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,35.1,446.1,1,28,58,0.0,3104,1,Fresno,0,0,Cable,36.878709,-119.7645,0,36.50400000000001,0,0,Offer D,45087,0,0,0,1,13,1,259.0,0.0,0.0,446.1,1,0,93720
5800,0,0,0,0,17,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),80.05,1345.65,0,62,29,44.96,3443,0,Fresno,1,0,Fiber Optic,36.732694,-119.783786,0,80.05,0,0,Offer D,6848,0,0,0,0,17,2,0.0,764.32,0.0,1345.65,0,1,93721
5801,1,1,1,0,34,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.55,2425.4,0,66,16,2.07,5381,0,Fresno,0,1,Cable,36.78979,-119.92989399999999,1,75.55,0,1,None,60889,0,0,1,0,34,0,388.0,70.38,0.0,2425.4,0,0,93722
5802,0,0,0,0,42,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,49.55,2077.95,0,40,23,8.71,3637,0,Fresno,0,0,DSL,36.623632,-119.741322,0,49.55,0,0,None,21010,0,0,0,0,42,0,0.0,365.82000000000005,0.0,2077.95,0,1,93725
5803,1,0,1,0,5,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,81.3,416.3,1,33,29,25.11,3819,1,Fresno,0,1,DSL,36.793601,-119.761131,1,84.552,0,0,Offer E,39148,0,2,0,0,5,6,121.0,125.55,0.0,416.3,0,0,93726
5804,0,0,1,1,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),23.9,1663.5,0,25,0,29.41,5471,0,Fresno,0,0,NA,36.751489,-119.68072,1,23.9,2,1,Offer A,54701,0,0,1,0,71,0,0.0,2088.11,0.0,1663.5,1,0,93727
5805,1,1,1,0,19,1,0,DSL,1,0,1,0,Month-to-month,0,Bank transfer (automatic),66.4,1286.05,0,71,26,30.44,4533,0,Fresno,1,1,Fiber Optic,36.757345,-119.818274,1,66.4,0,1,None,16346,0,0,1,0,19,0,0.0,578.36,0.0,1286.05,0,1,93728
5806,0,0,0,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.6,35.85,1,31,0,29.81,2843,1,Salinas,0,0,NA,36.64152,-121.622188,0,19.6,5,0,None,35739,0,1,0,0,2,3,0.0,59.62,0.0,35.85,0,0,93901
5807,1,0,0,0,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),18.8,1094.35,0,45,0,19.69,6466,0,Salinas,0,1,NA,36.667794,-121.60130600000001,0,18.8,0,0,None,58548,0,0,0,0,57,1,0.0,1122.3300000000004,0.0,1094.35,0,0,93905
5808,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,108.4,7719.5,0,29,59,10.68,4394,0,Salinas,1,1,Cable,36.722898,-121.633648,1,108.4,0,8,Offer A,53946,1,0,1,1,72,0,4555.0,768.96,0.0,7719.5,1,0,93906
5809,0,0,0,0,6,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Mailed check,85.95,514.6,0,28,51,40.64,3291,0,Salinas,0,0,DSL,36.77462,-121.66471399999999,0,85.95,0,0,None,22292,0,0,0,1,6,1,262.0,243.84,0.0,514.6,1,0,93907
5810,0,0,1,1,17,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.45,1451.6,1,29,29,47.76,3670,1,Salinas,0,0,Fiber Optic,36.624338,-121.615669,1,88.86800000000002,0,1,None,13027,0,1,1,1,17,4,0.0,811.92,0.0,1451.6,1,1,93908
5811,1,0,1,0,61,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),80.9,4932.5,0,29,51,23.31,4161,0,Escondido,1,1,Cable,33.141265000000004,-116.967221,1,80.9,0,1,None,48690,0,0,1,1,61,1,0.0,1421.91,0.0,4932.5,1,1,92027
5812,1,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,71.0,71,1,57,21,18.84,4207,1,Carmel By The Sea,0,1,Fiber Optic,36.554618,-121.92223899999999,1,73.84,0,1,Offer E,2966,0,0,1,0,1,2,0.0,18.84,0.0,71.0,0,0,93921
5813,1,0,1,1,48,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),111.8,5443.65,0,49,18,12.57,3922,0,Carmel,1,1,Fiber Optic,36.460611,-121.852507,1,111.8,2,10,None,13121,1,0,1,1,48,0,97.99,603.36,0.0,5443.65,0,1,93923
5814,1,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.6,330.25,0,36,0,33.44,5667,0,Carmel Valley,0,1,NA,36.414611,-121.6386,0,20.6,0,0,Offer D,6691,0,0,0,0,16,0,0.0,535.04,0.0,330.25,0,0,93924
5815,1,1,0,0,9,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.05,746.5,1,68,7,12.18,5095,1,Chualar,0,1,Cable,36.596271,-121.442274,0,88.45200000000001,0,0,Offer E,1140,0,0,0,0,9,7,0.0,109.62,0.0,746.5,0,1,93925
5816,0,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,44.6,122.7,0,62,27,15.59,3122,0,Gonzales,0,0,DSL,36.52588,-121.39671899999999,0,44.6,0,0,None,9023,0,0,0,0,3,2,33.0,46.77,0.0,122.7,0,0,93926
5817,1,0,0,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.4,44.4,1,29,57,7.14,4067,1,Greenfield,0,1,Fiber Optic,36.248708,-121.38661699999999,0,46.176,3,0,Offer E,14204,0,0,0,1,1,2,0.0,7.14,0.0,44.4,1,0,93927
5818,1,0,0,0,65,1,1,Fiber optic,0,1,1,1,Two year,0,Credit card (automatic),105.1,6631.85,0,47,30,27.75,5649,0,Jolon,1,1,Cable,35.930782,-121.189757,0,105.1,0,0,Offer B,254,0,0,0,1,65,0,198.96,1803.75,0.0,6631.85,0,1,93928
5819,0,0,1,1,70,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),115.15,8250,0,45,53,11.36,4388,0,King City,1,0,Cable,36.220760999999996,-120.980777,1,115.15,3,3,Offer A,14477,1,0,1,1,70,1,4372.0,795.1999999999998,0.0,8250.0,0,0,93930
5820,1,0,1,0,60,1,0,DSL,1,0,1,0,One year,1,Mailed check,59.8,3561.15,0,39,16,15.24,5488,0,Lockwood,0,1,Fiber Optic,35.989792,-121.05593300000001,1,59.8,0,6,Offer B,538,0,0,1,0,60,1,0.0,914.4,0.0,3561.15,0,1,93932
5821,0,0,1,0,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Electronic check,26.3,1763.55,0,23,0,22.08,5418,0,Marina,0,0,NA,36.689582,-121.758398,1,26.3,0,7,Offer A,21759,0,0,1,0,69,0,0.0,1523.52,0.0,1763.55,1,0,93933
5822,0,1,0,0,35,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.55,2419,0,65,30,16.91,5873,0,Monterey,0,0,DSL,36.362741,-121.869685,0,70.55,0,0,None,32857,0,0,0,0,35,0,0.0,591.85,0.0,2419.0,0,1,93940
5823,0,0,0,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.05,470.2,0,43,0,33.92,5555,0,Pacific Grove,0,0,NA,36.618337,-121.92641699999999,0,20.05,0,0,Offer D,15449,0,1,0,0,22,1,0.0,746.24,0.0,470.2,0,0,93950
5824,1,0,1,1,66,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),79.85,5234.95,0,25,59,35.01,6236,0,Pebble Beach,1,1,Fiber Optic,36.587497,-121.94481499999999,1,79.85,1,8,Offer A,4602,0,0,1,1,66,1,3089.0,2310.66,0.0,5234.95,1,0,93953
5825,1,1,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,70.3,1,80,30,39.1,4962,1,San Lucas,0,1,DSL,36.125529,-120.864443,1,73.112,0,0,Offer E,521,0,1,0,0,1,2,0.0,39.1,0.0,70.3,0,0,93954
5826,0,0,1,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),79.35,79.35,1,30,57,23.63,3492,1,Seaside,0,0,DSL,36.625114,-121.82356499999999,1,82.524,0,2,Offer E,38244,0,0,1,0,1,6,0.0,23.63,0.0,79.35,0,0,93955
5827,1,0,1,1,34,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),90.05,3097,0,61,57,20.05,4648,0,Soledad,1,1,Fiber Optic,36.414215999999996,-121.360597,1,90.05,3,10,Offer C,13003,0,0,1,1,34,2,1765.0,681.7,0.0,3097.0,0,0,93960
5828,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.45,1709.1,0,36,0,20.56,5335,0,Spreckels,0,0,NA,36.624641,-121.647195,1,24.45,1,4,Offer A,407,0,0,1,0,72,2,0.0,1480.32,0.0,1709.1,0,0,93962
5829,1,0,1,1,31,0,No phone service,DSL,1,0,1,1,One year,0,Electronic check,59.95,1848.8,0,64,25,0.0,4337,0,Belmont,1,1,Cable,37.509366,-122.306132,1,59.95,2,7,Offer C,25566,1,0,1,1,31,0,46.22,0.0,0.0,1848.8,0,1,94002
5830,1,0,0,1,30,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),25.35,723.3,0,61,0,4.27,5915,0,Brisbane,0,1,NA,37.684694,-122.40711999999999,0,25.35,2,0,Offer C,3635,0,0,0,0,30,1,0.0,128.1,0.0,723.3,0,0,94005
5831,0,0,0,0,9,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),90.8,809.75,1,53,10,1.34,2578,1,Burlingame,0,0,DSL,37.57028,-122.365778,0,94.432,0,0,Offer E,40346,0,1,0,1,9,1,0.0,12.06,0.0,809.75,0,1,94010
5832,1,0,1,1,20,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.45,1470.95,1,47,9,16.49,4773,1,Daly City,0,1,Cable,37.691561,-122.445202,1,73.268,0,1,None,47453,0,2,1,0,20,4,132.0,329.7999999999999,0.0,1470.95,0,0,94014
5833,1,1,1,0,19,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),34.3,577.15,0,65,14,0.0,4615,0,Daly City,1,1,Cable,37.680844,-122.48131000000001,1,34.3,0,6,None,63337,0,0,1,0,19,0,8.08,0.0,0.0,577.15,0,1,94015
5834,0,0,1,0,65,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,105.05,6914.95,0,35,23,40.71,5313,0,Half Moon Bay,1,0,DSL,37.45567,-122.407992,1,105.05,0,3,Offer B,17929,0,0,1,1,65,0,0.0,2646.15,0.0,6914.95,0,1,94019
5835,0,0,1,1,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.3,602.9,0,49,0,11.6,4453,0,La Honda,0,0,NA,37.285677,-122.22416499999999,1,19.3,1,8,Offer C,1622,0,0,1,0,30,0,0.0,348.0,0.0,602.9,0,0,94020
5836,1,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.15,124.4,0,33,0,10.54,5322,0,Loma Mar,0,1,NA,37.266388,-122.26308,0,19.15,0,0,None,148,0,1,0,0,6,1,0.0,63.24,0.0,124.4,0,0,94021
5837,0,0,0,0,2,0,No phone service,DSL,0,1,1,1,Month-to-month,0,Electronic check,51.4,96.8,0,53,21,0.0,2580,0,Los Altos,0,0,Fiber Optic,37.349546000000004,-122.13435600000001,0,51.4,0,0,None,18486,0,0,0,1,2,2,0.0,0.0,0.0,96.8,0,1,94022
5838,1,0,1,1,53,1,1,DSL,1,0,0,1,Month-to-month,0,Electronic check,71.85,3827.9,0,61,26,27.56,4903,0,Los Altos,0,1,DSL,37.352911,-122.093002,1,71.85,3,0,Offer B,21496,1,0,0,1,53,1,0.0,1460.6799999999996,0.0,3827.9,0,1,94024
5839,1,1,1,0,7,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.4,533.05,0,80,21,21.37,3533,0,Menlo Park,0,1,Fiber Optic,37.449551,-122.18376200000002,1,75.4,0,2,None,39062,0,0,1,0,7,2,0.0,149.59,0.0,533.05,0,1,94025
5840,0,0,1,1,61,1,0,DSL,1,0,0,0,One year,1,Bank transfer (automatic),49.7,2961.4,0,34,11,42.85,4577,0,Atherton,0,0,Fiber Optic,37.454924,-122.20316799999999,1,49.7,2,2,Offer B,6876,0,0,1,0,61,1,32.58,2613.85,0.0,2961.4,0,1,94027
5841,1,1,0,0,70,0,No phone service,DSL,0,0,1,1,One year,1,Electronic check,45.25,3264.45,1,79,22,0.0,5824,1,Portola Valley,0,1,DSL,37.369709,-122.21584399999999,0,47.06,0,0,None,6601,0,1,0,0,70,4,718.0,0.0,0.0,3264.45,0,0,94028
5842,0,0,0,0,13,1,1,DSL,1,0,1,1,Month-to-month,1,Electronic check,78.75,995.35,0,34,23,38.4,5631,0,Millbrae,1,0,Cable,37.601248,-122.403099,0,78.75,0,0,Offer D,20350,0,0,0,1,13,1,22.89,499.2,0.0,995.35,0,1,94030
5843,1,1,1,0,35,1,1,Fiber optic,0,0,0,0,One year,1,Bank transfer (automatic),81.6,2815.25,0,76,28,4.16,2300,0,Montara,1,1,DSL,37.540582,-122.50959399999999,1,81.6,0,2,None,2346,0,0,1,0,35,0,0.0,145.6,0.0,2815.25,0,1,94037
5844,0,0,1,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),70.4,154.8,0,61,14,7.49,5748,0,Moss Beach,0,0,DSL,37.515556,-122.502311,1,70.4,0,9,None,3064,0,0,1,0,2,0,22.0,14.98,0.0,154.8,0,0,94038
5845,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.8,246.3,1,63,25,5.2,5475,1,Mountain View,0,0,Fiber Optic,37.380662,-122.086022,0,78.832,0,0,Offer E,32143,0,1,0,0,3,3,62.0,15.6,0.0,246.3,0,0,94040
5846,0,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,76.1,257.6,0,50,17,14.35,2650,0,Mountain View,0,0,Fiber Optic,37.388349,-122.075299,0,76.1,0,0,None,13483,0,0,0,0,3,0,0.0,43.05,0.0,257.6,0,1,94041
5847,0,0,0,0,62,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),94.0,5757.2,0,42,26,32.29,4778,0,Mountain View,0,0,DSL,37.419725,-122.062947,0,94.0,0,0,Offer B,27822,0,0,0,1,62,0,149.69,2001.98,0.0,5757.2,0,1,94043
5848,1,0,1,1,72,1,1,Fiber optic,1,1,0,1,Two year,0,Credit card (automatic),103.95,7517.7,0,26,30,45.93,4495,0,Pacifica,1,1,Fiber Optic,37.573633,-122.45516699999999,1,103.95,2,1,Offer A,38885,1,1,1,1,72,3,2255.0,3306.96,0.0,7517.7,1,0,94044
5849,1,0,1,0,63,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.95,1234.8,0,56,0,38.36,5151,0,Pescadero,0,1,NA,37.22565,-122.297533,1,19.95,0,2,Offer B,2055,0,0,1,0,63,1,0.0,2416.68,0.0,1234.8,0,0,94060
5850,1,1,0,0,20,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),71.3,1389.2,1,78,24,5.71,3684,1,Redwood City,0,1,Fiber Optic,37.461251000000004,-122.23541399999999,0,74.152,0,0,Offer D,35737,0,0,0,0,20,2,333.0,114.2,0.0,1389.2,0,0,94061
5851,0,1,0,0,35,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),110.8,3836.3,0,74,22,32.92,2125,0,Redwood City,1,0,Fiber Optic,37.410567,-122.297152,0,110.8,0,0,None,25569,1,0,0,1,35,0,0.0,1152.2,0.0,3836.3,0,1,94062
5852,1,1,1,0,21,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.1,1474.75,1,76,20,19.74,3853,1,Redwood City,0,1,DSL,37.499411,-122.19631799999999,1,71.86399999999998,0,1,Offer D,32368,0,0,1,0,21,6,0.0,414.54,0.0,1474.75,0,1,94063
5853,1,0,1,0,62,1,1,Fiber optic,1,1,0,1,One year,0,Electronic check,96.1,6001.45,0,19,41,30.51,6139,0,Redwood City,0,1,Fiber Optic,37.527497,-122.23094099999999,1,96.1,0,4,Offer B,10658,0,0,1,1,62,1,246.06,1891.62,0.0,6001.45,1,1,94065
5854,0,0,0,0,15,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,48.8,720.1,0,34,18,26.54,2577,0,San Bruno,0,0,Fiber Optic,37.624435999999996,-122.43066100000001,0,48.8,0,0,Offer D,39566,0,0,0,0,15,1,130.0,398.1,0.0,720.1,0,0,94066
5855,0,0,0,0,55,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),50.55,2832.75,0,38,17,3.62,6250,0,San Carlos,0,0,DSL,37.497915,-122.26736100000001,0,50.55,0,0,Offer B,28098,0,0,0,0,55,1,0.0,199.1,0.0,2832.75,0,1,94070
5856,0,0,0,0,11,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.65,472.25,0,59,3,29.16,4492,0,San Gregorio,0,0,Cable,37.331762,-122.341444,0,44.65,0,0,Offer D,291,0,0,0,0,11,0,0.0,320.76,0.0,472.25,0,1,94074
5857,0,0,1,1,17,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,88.25,1460.65,1,31,10,17.91,4041,1,South San Francisco,1,0,DSL,37.654436,-122.426468,1,91.78,0,7,None,60599,0,0,1,0,17,2,146.0,304.47,0.0,1460.65,0,0,94080
5858,0,0,0,0,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),19.45,1336.35,0,24,0,25.91,4559,0,Sunnyvale,0,0,NA,37.378541,-122.02045600000001,0,19.45,0,0,Offer B,64010,0,2,0,0,61,2,0.0,1580.51,0.0,1336.35,1,0,94086
5859,0,0,1,0,71,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.3,6388.65,0,38,27,19.9,4658,0,Sunnyvale,1,0,Cable,37.3511,-122.03731100000002,1,89.3,0,7,Offer A,50070,1,0,1,1,71,0,0.0,1412.9,0.0,6388.65,0,1,94087
5860,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),70.0,153.05,1,31,11,37.76,2928,1,Sunnyvale,0,0,Fiber Optic,37.421633,-122.00961299999999,0,72.8,0,0,Offer E,16985,0,0,0,0,2,2,17.0,75.52,0.0,153.05,0,0,94089
5861,1,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.25,677.9,0,33,0,4.24,2682,0,San Francisco,0,1,NA,37.7795,-122.419233,0,19.25,0,0,Offer C,28998,0,0,0,0,35,0,0.0,148.4,0.0,677.9,0,0,94102
5862,0,0,0,0,17,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),70.5,1165.6,0,53,16,41.78,3650,0,San Francisco,0,0,DSL,37.773146999999994,-122.41128700000002,0,70.5,0,0,Offer D,23036,0,0,0,0,17,1,0.0,710.26,0.0,1165.6,0,1,94103
5863,0,0,0,0,21,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,97.35,2119.5,1,63,11,9.06,4321,1,San Francisco,0,0,Cable,37.791222,-122.40224099999999,0,101.244,0,0,None,384,0,0,0,1,21,3,233.0,190.26,0.0,2119.5,0,0,94104
5864,0,0,1,0,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.65,921.55,0,21,0,45.9,4159,0,San Francisco,0,0,NA,37.789168,-122.395009,1,19.65,0,1,Offer B,2066,0,0,1,0,47,1,0.0,2157.3,0.0,921.55,1,0,94105
5865,0,0,1,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.85,72,0,35,0,11.77,5867,0,San Francisco,0,0,NA,37.768881,-122.395521,1,20.85,0,9,None,17372,0,2,1,0,3,1,0.0,35.31,0.0,72.0,0,0,94107
5866,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.65,68.35,0,46,0,35.59,4852,0,San Francisco,0,1,NA,37.791998,-122.408653,0,19.65,0,0,None,13723,0,0,0,0,3,0,0.0,106.77,0.0,68.35,0,0,94108
5867,1,1,1,0,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.35,847.25,0,74,0,1.89,4975,0,San Francisco,0,1,NA,37.794487,-122.42227,1,19.35,0,4,None,56330,0,0,1,0,44,2,0.0,83.16,0.0,847.25,0,0,94109
5868,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.0,44,0,51,26,26.15,4138,0,San Francisco,0,0,Fiber Optic,37.750021000000004,-122.415201,0,44.0,0,0,None,74641,0,1,0,0,1,1,0.0,26.15,0.0,44.0,0,1,94110
5869,0,0,1,1,44,1,1,Fiber optic,0,1,0,1,One year,0,Electronic check,94.4,4295.35,0,40,27,24.71,5019,0,San Francisco,1,0,DSL,37.801776000000004,-122.402293,1,94.4,2,4,Offer B,3337,0,0,1,1,44,0,0.0,1087.24,0.0,4295.35,0,1,94111
5870,1,0,1,1,5,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Bank transfer (automatic),25.9,135,1,34,0,40.05,2102,1,San Francisco,0,1,NA,37.720498,-122.443119,1,25.9,1,1,Offer E,73117,0,0,1,0,5,3,0.0,200.25,0.0,135.0,0,0,94112
5871,1,0,0,0,24,1,1,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),55.65,1400.55,1,43,6,8.99,4126,1,San Francisco,0,1,DSL,37.758084999999994,-122.43480100000001,0,57.876000000000005,0,0,None,30587,0,2,0,0,24,2,84.0,215.76,0.0,1400.55,0,0,94114
5872,0,0,0,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.65,69.65,1,52,9,49.24,2418,1,San Francisco,0,0,Cable,37.786031,-122.437301,0,72.436,0,0,Offer E,33122,0,0,0,0,1,2,0.0,49.24,0.0,69.65,0,1,94115
5873,0,0,0,0,18,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,75.4,1380.4,0,44,22,15.01,4792,0,San Francisco,0,0,DSL,37.744409999999995,-122.486764,0,75.4,0,0,Offer D,42959,0,0,0,0,18,1,0.0,270.18,0.0,1380.4,0,1,94116
5874,0,0,0,0,10,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.6,1060.2,1,41,3,45.21,4001,1,San Francisco,1,0,Fiber Optic,37.770533,-122.445121,0,104.624,0,0,None,38756,0,2,0,1,10,2,32.0,452.1,0.0,1060.2,0,0,94117
5875,0,0,1,0,65,1,0,DSL,1,1,0,1,Two year,0,Bank transfer (automatic),71.0,4386.2,0,25,51,1.29,6308,0,San Francisco,1,0,DSL,37.781304,-122.461522,1,71.0,0,1,Offer B,38955,0,0,1,1,65,0,0.0,83.85000000000002,0.0,4386.2,1,1,94118
5876,0,1,0,0,1,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,86.0,86,1,65,24,28.82,5359,1,San Francisco,0,0,DSL,37.776718,-122.49578100000001,0,89.44,0,0,Offer E,42476,0,0,0,1,1,4,0.0,28.82,0.0,86.0,0,0,94121
5877,0,0,0,0,53,1,1,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),106.95,5785.5,1,44,4,29.8,5550,1,San Francisco,1,0,Cable,37.760412,-122.48496599999999,0,111.228,0,0,None,55504,0,1,0,1,53,1,231.0,1579.4,0.0,5785.5,0,0,94122
5878,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,21.2,52.05,0,40,0,12.05,2088,0,San Francisco,0,1,NA,37.800253999999995,-122.436975,0,21.2,0,0,None,22920,0,0,0,0,3,0,0.0,36.15000000000001,0.0,52.05,0,0,94123
5879,1,0,1,0,33,1,0,DSL,1,1,0,0,Two year,1,Mailed check,61.05,2018.4,0,19,52,15.89,3215,0,San Francisco,0,1,Cable,37.731505,-122.38453200000001,1,61.05,0,3,Offer C,33177,1,0,1,0,33,0,1050.0,524.37,0.0,2018.4,1,0,94124
5880,1,0,0,0,3,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Electronic check,29.6,79.45,1,46,3,0.0,2734,1,San Francisco,0,1,DSL,37.736534999999996,-122.45732,0,30.784,0,0,Offer E,20643,0,1,0,0,3,3,2.0,0.0,0.0,79.45,0,0,94127
5881,0,0,0,0,34,1,0,DSL,1,0,1,1,One year,1,Bank transfer (automatic),79.95,2727.3,0,40,23,5.32,3570,0,San Francisco,1,0,DSL,37.797526,-122.46453100000001,0,79.95,0,0,Offer C,2240,1,0,0,1,34,0,627.0,180.88,0.0,2727.3,0,0,94129
5882,0,0,1,1,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.7,263.65,0,40,0,15.33,2966,0,San Francisco,0,0,NA,37.820894,-122.369725,1,19.7,1,8,Offer D,1458,0,0,1,0,14,2,0.0,214.62,0.0,263.65,0,0,94130
5883,0,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.3,275.4,0,27,0,22.01,5332,0,San Francisco,0,0,NA,37.746699,-122.44283300000001,0,20.3,0,0,Offer D,27906,0,0,0,0,13,0,0.0,286.13,0.0,275.4,1,0,94131
5884,1,1,1,0,46,0,No phone service,DSL,0,1,1,1,One year,1,Bank transfer (automatic),59.9,2816.65,1,80,16,0.0,4011,1,San Francisco,1,1,DSL,37.722302,-122.491129,1,62.29600000000001,0,1,None,26297,1,0,1,0,46,2,451.0,0.0,0.0,2816.65,0,0,94132
5885,1,0,1,1,23,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,24.35,538.5,0,22,0,48.02,4031,0,San Francisco,0,1,NA,37.802071000000005,-122.411004,1,24.35,3,1,None,26831,0,0,1,0,23,0,0.0,1104.46,0.0,538.5,1,0,94133
5886,0,0,1,1,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,948.9,0,33,0,41.54,3843,0,San Francisco,0,0,NA,37.721052,-122.413573,1,19.75,3,10,Offer B,40137,0,0,1,0,47,1,0.0,1952.38,0.0,948.9,0,0,94134
5887,1,0,0,1,17,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,50.3,846.8,0,35,53,45.61,3202,0,Palo Alto,0,1,DSL,37.444314,-122.149996,0,50.3,3,0,None,16198,0,0,0,0,17,0,0.0,775.37,0.0,846.8,0,1,94301
5888,0,0,1,1,49,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.6,4783.5,1,53,10,49.63,5732,1,Palo Alto,0,0,Cable,37.458090000000006,-122.115398,1,99.424,0,2,None,45499,0,0,1,1,49,3,478.0,2431.870000000001,0.0,4783.5,0,0,94303
5889,1,1,1,0,59,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,50.25,2997.45,0,65,23,0.0,5546,0,Palo Alto,0,1,Cable,37.386978000000006,-122.177746,1,50.25,0,4,None,1723,0,0,1,1,59,1,689.0,0.0,0.0,2997.45,0,0,94304
5890,0,0,0,0,69,1,1,DSL,1,0,1,1,Two year,1,Credit card (automatic),85.35,5897.4,0,42,28,18.47,6499,0,Stanford,1,0,Fiber Optic,37.424341999999996,-122.165641,0,85.35,0,0,Offer A,13386,1,0,0,1,69,0,165.13,1274.4299999999996,0.0,5897.4,0,1,94305
5891,1,0,0,0,11,0,No phone service,DSL,0,0,1,0,One year,1,Electronic check,41.6,470.6,1,39,6,0.0,3119,1,Palo Alto,1,1,Fiber Optic,37.416159,-122.13133700000002,0,43.263999999999996,0,0,None,24492,0,1,0,0,11,3,0.0,0.0,0.0,470.6,0,1,94306
5892,1,0,0,0,10,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,51.65,524.5,0,38,23,49.04,4292,0,San Mateo,0,1,Fiber Optic,37.590421,-122.306467,0,51.65,0,0,None,32488,0,2,0,0,10,1,0.0,490.4,0.0,524.5,0,1,94401
5893,1,0,1,1,12,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.0,269.65,0,56,0,26.17,3705,0,San Mateo,0,1,NA,37.556634,-122.317723,1,24.0,1,0,None,23393,0,0,0,0,12,0,0.0,314.04,0.0,269.65,0,0,94402
5894,1,0,0,0,45,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),100.85,4740,1,34,3,14.12,4898,1,San Mateo,0,1,Cable,37.538309000000005,-122.305109,0,104.884,0,0,Offer B,37926,0,0,0,1,45,1,142.0,635.4,0.0,4740.0,0,0,94403
5895,0,0,1,1,39,1,0,DSL,0,0,1,0,Month-to-month,1,Mailed check,59.85,2341.5,0,32,23,48.14,3900,0,San Mateo,1,0,DSL,37.556094,-122.27243700000001,1,59.85,2,4,Offer C,31882,0,0,1,0,39,0,0.0,1877.46,0.0,2341.5,0,1,94404
5896,1,1,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.45,1789.65,0,80,0,37.25,5341,0,Alameda,0,1,NA,37.774633,-122.27443400000001,1,25.45,0,3,Offer A,58555,0,1,1,0,71,2,0.0,2644.75,0.0,1789.65,0,0,94501
5897,1,0,1,1,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),23.9,1626.4,0,39,0,18.99,5574,0,Alameda,0,1,NA,37.724817,-122.22436299999998,1,23.9,1,9,Offer A,13996,0,0,1,0,71,1,0.0,1348.29,0.0,1626.4,0,0,94502
5898,0,0,1,1,33,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),24.15,800.3,0,22,0,1.71,4501,0,Danville,0,0,NA,37.791481,-121.903253,1,24.15,1,3,Offer C,19777,0,0,1,0,33,1,0.0,56.43,0.0,800.3,1,0,94506
5899,1,1,0,0,67,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,75.7,5060.85,0,75,19,39.89,5823,0,Alamo,0,1,Fiber Optic,37.855717,-121.994813,0,75.7,0,0,Offer A,15187,0,0,0,0,67,0,0.0,2672.63,0.0,5060.85,0,1,94507
5900,1,0,1,1,37,0,No phone service,DSL,1,1,0,0,Month-to-month,0,Bank transfer (automatic),40.2,1448.8,1,52,25,0.0,3627,1,Angwin,1,1,Cable,38.542448,-122.419923,1,41.80800000000001,1,1,None,3641,0,0,1,0,37,2,362.0,0.0,0.0,1448.8,0,0,94508
5901,1,0,1,1,49,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,84.5,4254.85,1,55,22,39.6,4639,1,Antioch,0,1,Cable,37.980057,-121.801599,1,87.88000000000002,0,1,Offer B,90891,0,0,1,0,49,2,936.0,1940.4,0.0,4254.85,0,0,94509
5902,0,0,1,0,9,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,50.85,466.6,0,19,76,12.59,4623,0,Benicia,0,0,Fiber Optic,38.113533000000004,-122.11926000000001,1,50.85,0,4,None,25578,0,0,1,0,9,2,355.0,113.31,0.0,466.6,1,0,94510
5903,1,0,1,0,52,1,1,Fiber optic,1,0,0,0,Two year,1,Credit card (automatic),91.6,4627.8,0,61,3,18.02,6069,0,Bethel Island,1,1,DSL,38.050558,-121.646924,1,91.6,0,3,Offer B,2379,1,0,1,0,52,1,0.0,937.04,0.0,4627.8,0,1,94511
5904,0,0,0,0,70,1,1,Fiber optic,0,1,1,1,One year,0,Electronic check,98.9,6838.6,0,25,59,8.39,5980,0,Birds Landing,0,0,DSL,38.140719,-121.838298,0,98.9,0,0,Offer A,138,0,0,0,1,70,0,4035.0,587.3000000000002,0.0,6838.6,1,0,94512
5905,1,0,0,0,1,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,85.0,85,0,60,2,15.2,5754,0,Brentwood,0,1,Fiber Optic,37.908242,-121.682472,0,85.0,0,0,None,26577,0,0,0,1,1,0,0.0,15.2,0.0,85.0,0,1,94513
5906,0,1,0,0,14,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,78.95,1101.85,1,65,7,16.36,5203,1,Byron,0,0,Fiber Optic,37.83323,-121.60146100000001,0,82.10799999999999,0,0,Offer D,10153,0,0,0,0,14,2,77.0,229.04,0.0,1101.85,0,0,94514
5907,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,44.3,44.3,0,54,9,42.95,4427,0,Calistoga,0,1,Cable,38.629618,-122.593216,0,44.3,0,0,Offer E,7384,0,0,0,0,1,0,0.0,42.95,0.0,44.3,0,0,94515
5908,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.2,20.2,1,45,0,11.25,5418,1,Clayton,0,1,NA,37.881842,-121.84811100000002,0,20.2,0,0,Offer E,14239,0,0,0,0,1,0,0.0,11.25,0.0,20.2,0,0,94517
5909,0,0,0,0,52,1,1,Fiber optic,0,1,0,0,One year,1,Mailed check,80.2,4297.6,0,43,14,42.9,5597,0,Concord,0,0,Fiber Optic,37.950247999999995,-122.02245500000001,0,80.2,0,0,Offer B,27394,0,0,0,0,52,2,0.0,2230.8,0.0,4297.6,0,1,94518
5910,1,0,0,0,6,1,0,DSL,0,0,1,0,Month-to-month,0,Mailed check,60.9,414.1,0,29,71,45.67,2191,0,Concord,1,1,Fiber Optic,37.990118,-122.012188,0,60.9,0,0,Offer E,18650,0,0,0,0,6,0,294.0,274.02,0.0,414.1,1,0,94519
5911,1,0,1,0,7,0,No phone service,DSL,1,1,0,0,Month-to-month,0,Mailed check,34.2,256.6,0,47,17,0.0,5100,0,Concord,0,1,Cable,38.013825,-122.039144,1,34.2,0,3,Offer E,36186,0,0,1,0,7,0,0.0,0.0,0.0,256.6,0,1,94520
5912,0,1,0,0,47,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),85.2,3969.35,1,78,13,16.83,4661,1,Concord,1,0,DSL,37.971421,-121.97150400000001,0,88.60799999999999,0,0,None,39888,0,1,0,0,47,1,516.0,791.0099999999999,0.0,3969.35,0,0,94521
5913,0,0,0,0,26,1,0,Fiber optic,1,0,0,0,One year,1,Credit card (automatic),87.15,2274.1,0,19,41,45.09,5689,0,Pleasant Hill,1,0,DSL,37.953379999999996,-122.07688600000002,0,87.15,0,0,Offer C,32685,1,0,0,0,26,1,0.0,1172.34,0.0,2274.1,1,1,94523
5914,1,0,1,1,25,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,54.3,1296.8,0,34,22,37.97,3971,0,Crockett,0,1,Fiber Optic,38.049292,-122.22841499999998,1,54.3,1,6,Offer C,3193,1,0,1,0,25,2,285.0,949.25,0.0,1296.8,0,0,94525
5915,1,0,0,0,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.1,1268.85,0,19,0,42.49,4535,0,Danville,0,1,NA,37.815459000000004,-121.977203,0,19.1,0,0,Offer A,32873,0,0,0,0,69,0,0.0,2931.81,0.0,1268.85,1,0,94526
5916,0,0,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),112.75,8192.6,0,30,42,35.24,4927,0,El Cerrito,1,0,DSL,37.924838,-122.28914499999999,0,112.75,0,0,Offer A,23141,1,0,0,1,72,0,0.0,2537.28,0.0,8192.6,0,1,94530
5917,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.95,59.25,0,55,0,34.86,3172,0,Fairfield,0,1,NA,38.287136,-122.02711000000001,0,19.95,0,0,None,77683,0,0,0,0,4,0,0.0,139.44,0.0,59.25,0,0,94533
5918,1,0,1,1,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.5,1147.85,0,35,0,18.75,5293,0,Travis Afb,0,1,NA,38.265899,-121.93946100000001,1,19.5,2,10,Offer B,9978,0,2,1,0,59,2,0.0,1106.25,0.0,1147.85,0,0,94535
5919,1,0,0,0,67,1,0,DSL,1,0,0,1,Two year,0,Bank transfer (automatic),65.55,4361.55,0,29,41,49.74,6035,0,Fremont,1,1,Fiber Optic,37.572272999999996,-121.964583,0,65.55,0,0,Offer A,66543,0,0,0,1,67,2,1788.0,3332.58,0.0,4361.55,1,0,94536
5920,0,1,0,0,26,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,78.8,2006.1,0,70,15,19.21,4509,0,Fremont,0,0,Fiber Optic,37.505767999999996,-121.96247199999999,0,78.8,0,0,None,56126,0,0,0,1,26,1,0.0,499.46,0.0,2006.1,0,1,94538
5921,0,0,0,0,27,1,0,DSL,0,1,1,1,One year,0,Mailed check,78.2,2078.95,0,20,59,48.91,2297,0,Fremont,1,0,DSL,37.516791,-121.89911699999999,0,78.2,0,0,Offer C,46917,1,0,0,1,27,0,1227.0,1320.57,0.0,2078.95,1,0,94539
5922,1,0,1,1,72,1,1,Fiber optic,1,0,1,1,Two year,0,Bank transfer (automatic),105.25,7609.75,0,41,14,36.05,4427,0,Hayward,1,1,Cable,37.674002,-122.076796,1,105.25,2,5,Offer A,60274,0,0,1,1,72,1,1065.0,2595.6,0.0,7609.75,0,0,94541
5923,0,0,0,0,6,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.25,487.05,0,60,10,35.88,4430,0,Hayward,1,0,DSL,37.656695,-122.04836100000001,0,89.25,0,0,Offer E,11147,1,0,0,1,6,0,4.87,215.28000000000003,0.0,487.05,0,1,94542
5924,1,0,1,1,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.65,1218.45,0,55,0,11.15,6403,0,Hayward,0,1,NA,37.639215,-122.037554,1,20.65,2,9,Offer B,72993,0,0,1,0,62,1,0.0,691.3000000000002,0.0,1218.45,0,0,94544
5925,1,0,0,0,20,1,1,DSL,0,1,1,0,One year,1,Electronic check,68.7,1416.2,0,23,52,32.5,2989,0,Hayward,0,1,DSL,37.62984,-122.120843,0,68.7,0,0,None,27311,1,0,0,0,20,0,0.0,650.0,0.0,1416.2,1,1,94545
5926,1,0,0,0,6,1,0,DSL,1,0,1,1,Month-to-month,0,Credit card (automatic),78.65,483.3,0,44,7,46.59,2724,0,Castro Valley,1,1,DSL,37.708327000000004,-122.083473,0,78.65,0,0,Offer E,41698,1,0,0,1,6,1,0.0,279.54,0.0,483.3,0,1,94546
5927,1,0,0,0,51,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.75,1234.6,0,63,0,18.07,5080,0,Hercules,0,1,NA,37.991259,-122.214945,0,24.75,0,0,Offer B,22479,0,0,0,0,51,1,0.0,921.57,0.0,1234.6,0,0,94547
5928,0,0,1,1,61,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.75,1311.6,0,44,0,25.4,6108,0,Lafayette,0,0,NA,37.907777,-122.12716100000002,1,19.75,2,6,Offer B,23996,0,0,1,0,61,0,0.0,1549.4,0.0,1311.6,0,0,94549
5929,1,1,1,0,62,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,89.1,5618.3,0,68,3,4.76,4415,0,Livermore,1,1,Cable,37.571748,-121.65956200000001,1,89.1,0,4,None,75929,0,0,1,0,62,0,0.0,295.12,0.0,5618.3,0,1,94550
5930,0,0,0,0,72,1,1,Fiber optic,1,0,0,0,Two year,1,Bank transfer (automatic),84.7,6185.15,0,45,22,8.48,4520,0,Castro Valley,0,0,DSL,37.722727,-122.02157,0,84.7,0,0,Offer A,13212,1,0,0,0,72,1,0.0,610.5600000000002,0.0,6185.15,0,1,94552
5931,1,1,1,0,13,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,98.0,1237.85,1,78,4,27.82,3714,1,Martinez,1,1,DSL,38.014457,-122.11543200000001,1,101.92,0,1,Offer D,46677,0,0,1,0,13,0,50.0,361.66,0.0,1237.85,0,0,94553
5932,1,0,1,0,5,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.45,498.1,1,43,26,39.36,4580,1,Fremont,1,1,Cable,37.555473,-122.080312,1,98.228,0,1,None,33883,0,1,1,1,5,4,130.0,196.8,0.0,498.1,0,0,94555
5933,1,1,0,0,3,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.0,294.45,1,68,20,35.43,5960,1,Moraga,1,1,Cable,37.827946000000004,-122.10718500000002,0,109.2,0,0,Offer E,16510,0,1,0,0,3,5,59.0,106.29,0.0,294.45,0,0,94556
5934,0,1,1,0,26,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,93.85,2381.55,1,73,29,9.28,2591,1,Napa,1,0,Cable,38.489789,-122.27011,1,97.604,0,1,Offer C,63947,0,3,1,0,26,4,691.0,241.28,0.0,2381.55,0,0,94558
5935,1,1,0,0,13,1,0,DSL,0,1,1,0,Month-to-month,1,Electronic check,59.9,788.35,0,76,30,49.9,5254,0,Napa,0,1,Fiber Optic,38.232389000000005,-122.32494399999999,0,59.9,0,0,None,26894,0,0,0,0,13,0,0.0,648.6999999999998,0.0,788.35,0,1,94559
5936,0,0,1,1,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.95,756.4,0,26,0,49.9,3614,0,Newark,0,0,NA,37.504133,-122.032347,1,19.95,3,7,Offer C,42491,0,0,1,0,38,0,0.0,1896.2,0.0,756.4,1,0,94560
5937,0,1,1,0,8,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.0,613.4,1,75,24,46.05,4819,1,Oakley,0,0,Cable,37.999406,-121.686241,1,87.36,0,1,None,27607,0,1,1,0,8,6,0.0,368.4,0.0,613.4,0,1,94561
5938,1,1,1,1,34,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,108.9,3625.2,0,70,12,11.74,5151,0,Orinda,1,1,Fiber Optic,37.873915999999994,-122.20522,1,108.9,1,7,None,17964,1,0,1,1,34,1,0.0,399.16,0.0,3625.2,0,1,94563
5939,1,0,0,0,18,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,33.6,550.35,0,53,30,0.0,5388,0,Pinole,1,1,Cable,37.996462,-122.29371599999999,0,33.6,0,0,None,16717,0,0,0,0,18,0,165.0,0.0,0.0,550.35,0,0,94564
5940,1,0,1,1,56,1,0,Fiber optic,0,1,0,0,One year,1,Mailed check,85.85,4793.8,0,60,10,11.48,5058,0,Pittsburg,1,1,Fiber Optic,38.006046999999995,-121.91683400000001,1,85.85,1,4,None,78816,1,0,1,0,56,1,479.0,642.88,0.0,4793.8,0,0,94565
5941,0,0,0,0,36,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Bank transfer (automatic),34.85,1267.2,0,41,2,0.0,4452,0,Pleasanton,0,0,Fiber Optic,37.633361,-121.86239499999999,0,34.85,0,0,Offer C,36669,1,0,0,0,36,3,0.0,0.0,0.0,1267.2,0,1,94566
5942,0,0,1,0,9,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,48.75,442.2,1,51,11,0.0,4359,1,Pope Valley,1,0,Cable,38.672708,-122.40321899999999,1,50.7,0,1,None,494,0,0,1,1,9,2,49.0,0.0,0.0,442.2,0,0,94567
5943,1,0,0,0,1,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,84.85,84.85,1,25,45,36.07,3086,1,Dublin,1,1,DSL,37.713926,-121.928425,0,88.244,0,0,None,29636,0,1,0,1,1,2,0.0,36.07,0.0,84.85,1,0,94568
5944,1,0,0,0,12,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,56.65,654.85,1,42,11,7.97,3043,1,Port Costa,0,1,Cable,38.035707,-122.196821,0,58.916,0,0,None,173,1,2,0,0,12,4,0.0,95.64,0.0,654.85,0,1,94569
5945,0,1,1,1,57,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),95.3,5567.45,0,75,15,28.25,4912,0,Rio Vista,1,0,Fiber Optic,38.148862,-121.737696,1,95.3,1,8,None,5246,1,0,1,0,57,0,835.0,1610.25,0.0,5567.45,0,0,94571
5946,0,0,0,0,42,1,0,DSL,1,1,0,1,One year,0,Credit card (automatic),73.9,3160.55,1,22,58,5.75,2774,1,Rodeo,1,0,Fiber Optic,38.027218,-122.23463000000001,0,76.85600000000002,0,0,Offer B,8506,1,0,0,1,42,3,1833.0,241.5,0.0,3160.55,1,0,94572
5947,0,0,1,1,33,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.5,740.3,1,21,0,35.31,5194,1,Saint Helena,0,0,NA,38.581354,-122.296283,1,24.5,0,1,None,9423,0,0,1,0,33,0,0.0,1165.23,35.05,740.3,1,0,94574
5948,1,0,1,0,70,1,0,Fiber optic,1,1,0,0,Two year,0,Bank transfer (automatic),84.6,5706.2,0,45,21,1.07,5679,0,Deer Park,0,1,Fiber Optic,38.554383,-122.474773,1,84.6,0,3,Offer A,223,1,0,1,0,70,0,1198.0,74.9,0.0,5706.2,0,0,94576
5949,0,0,0,0,68,0,No phone service,DSL,0,1,0,1,Month-to-month,0,Electronic check,44.95,3085.35,0,53,13,0.0,5750,0,San Leandro,0,0,DSL,37.717196,-122.15933799999999,0,44.95,0,0,None,41871,1,0,0,1,68,1,401.0,0.0,0.0,3085.35,0,0,94577
5950,1,0,0,1,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,24.7,24.7,0,47,21,0.0,3518,0,San Leandro,0,1,DSL,37.704384000000005,-122.126703,0,24.7,3,0,None,36568,0,0,0,0,1,1,0.0,0.0,0.0,24.7,0,1,94578
5951,0,0,0,0,37,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Credit card (automatic),100.3,3541.4,0,26,82,45.06,4040,0,San Leandro,0,0,Cable,37.687264,-122.15728,0,100.3,0,0,None,19815,1,0,0,1,37,0,2904.0,1667.22,0.0,3541.4,1,0,94579
5952,0,0,0,1,4,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,25.45,84.2,0,20,0,38.97,2616,0,San Lorenzo,0,0,NA,37.676249,-122.132415,0,25.45,3,0,Offer E,26240,0,0,0,0,4,0,0.0,155.88,0.0,84.2,1,0,94580
5953,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,50.7,50.7,0,56,14,38.05,3007,0,San Ramon,0,1,Cable,37.766556,-121.97678400000001,0,50.7,0,0,Offer E,44078,0,0,0,0,1,1,0.0,38.05,0.0,50.7,0,0,94583
5954,1,0,0,0,20,0,No phone service,DSL,1,1,1,0,Month-to-month,1,Credit card (automatic),55.0,1165.55,0,45,20,0.0,4481,0,Suisun City,1,1,Fiber Optic,38.197907,-122.01725800000001,0,55.0,0,0,None,39279,1,0,0,0,20,3,23.31,0.0,0.0,1165.55,0,1,94585
5955,1,0,1,1,72,1,0,DSL,1,1,1,0,Two year,0,Bank transfer (automatic),68.4,4855.35,0,52,26,15.96,5504,0,Sunol,0,1,DSL,37.587494,-121.86285600000001,1,68.4,1,7,None,790,1,0,1,0,72,0,1262.0,1149.12,0.0,4855.35,0,0,94586
5956,0,0,0,0,31,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.9,2806.9,1,54,12,6.33,2031,1,Union City,1,0,DSL,37.59485,-122.051521,0,93.496,0,0,None,66472,0,3,0,1,31,3,337.0,196.23,41.18,2806.9,0,0,94587
5957,1,1,1,0,18,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,78.55,1422.65,1,66,20,4.98,3521,1,Pleasanton,0,1,Fiber Optic,37.685052,-121.91206100000001,1,81.692,0,1,Offer D,28568,0,2,1,0,18,1,285.0,89.64000000000001,0.0,1422.65,0,0,94588
5958,1,0,1,0,11,1,0,DSL,0,0,1,0,Month-to-month,1,Bank transfer (automatic),55.05,608.15,0,38,15,44.2,2762,0,Vallejo,0,1,Fiber Optic,38.161321,-122.271588,1,55.05,0,6,None,42209,0,0,1,0,11,1,91.0,486.2000000000001,0.0,608.15,0,0,94589
5959,0,0,1,1,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.8,641.35,0,35,0,12.51,2635,0,Vallejo,0,0,NA,38.104704999999996,-122.24738700000002,1,19.8,1,0,None,37218,0,0,0,0,33,1,0.0,412.83,0.0,641.35,0,0,94590
5960,0,1,0,0,62,1,1,Fiber optic,0,0,1,0,One year,0,Electronic check,84.45,4959.15,0,69,3,19.52,4166,0,Vallejo,0,0,DSL,38.105733,-122.18633799999999,0,84.45,0,0,None,51665,0,0,0,0,62,1,0.0,1210.24,0.0,4959.15,0,1,94591
5961,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,35.9,35.9,0,60,7,0.0,3929,0,Vallejo,1,0,Fiber Optic,38.093701,-122.27658899999999,0,35.9,0,0,Offer E,159,1,0,0,0,1,0,0.0,0.0,0.0,35.9,0,1,94592
5962,1,0,1,0,16,1,0,Fiber optic,1,1,0,0,Month-to-month,0,Bank transfer (automatic),80.75,1321.3,0,59,30,46.0,2942,0,Walnut Creek,0,1,DSL,37.862128000000006,-122.075197,1,80.75,0,8,None,18024,0,0,1,0,16,2,0.0,736.0,0.0,1321.3,0,1,94595
5963,1,0,1,1,22,1,1,DSL,0,0,1,1,One year,1,Mailed check,78.65,1663.75,0,64,11,36.15,3571,0,Walnut Creek,1,1,DSL,37.900662,-122.05278200000001,1,78.65,2,6,None,40917,1,0,1,1,22,1,183.0,795.3,0.0,1663.75,0,0,94596
5964,0,0,1,1,49,1,0,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),61.75,3024.15,0,35,28,35.29,5511,0,Walnut Creek,1,0,DSL,37.916647999999995,-122.00848300000001,1,61.75,1,6,None,26022,1,0,1,0,49,2,847.0,1729.21,0.0,3024.15,0,0,94598
5965,1,0,1,1,36,1,0,DSL,1,0,0,1,One year,1,Credit card (automatic),63.7,2188.5,0,36,14,47.45,2504,0,Yountville,1,1,Fiber Optic,38.421458,-122.365048,1,63.7,2,8,None,2873,0,1,1,1,36,1,306.0,1708.2,0.0,2188.5,0,0,94599
5966,1,0,1,0,42,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,99.45,4138.05,1,50,10,34.65,4624,1,Oakland,1,1,Cable,37.776523,-122.219268,1,103.428,0,1,Offer B,54876,1,2,1,1,42,1,414.0,1455.3,30.46,4138.05,0,0,94601
5967,1,1,0,0,4,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),25.2,102.5,1,73,21,0.0,4694,1,Oakland,0,1,Cable,37.803883,-122.208417,0,26.208000000000002,0,0,Offer E,28900,0,0,0,0,4,2,22.0,0.0,0.0,102.5,0,0,94602
5968,0,0,0,0,12,1,1,DSL,0,0,1,1,One year,0,Mailed check,74.05,872.65,1,57,24,42.58,4149,1,Oakland,0,0,DSL,37.739113,-122.175602,0,77.012,0,0,None,31392,1,0,0,1,12,2,0.0,510.96,48.61,872.65,0,1,94603
5969,0,0,0,0,31,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Electronic check,87.6,2724.25,0,56,20,40.92,5094,0,Oakland,1,0,DSL,37.758019,-122.138678,0,87.6,0,0,None,42854,1,0,0,0,31,2,0.0,1268.52,0.0,2724.25,0,1,94605
5970,1,0,1,0,5,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,89.15,413.25,0,33,28,15.74,2576,0,Oakland,0,1,Fiber Optic,37.792489,-122.24431399999999,1,89.15,0,8,Offer E,41876,0,0,1,1,5,1,0.0,78.7,0.0,413.25,0,1,94606
5971,1,0,1,1,66,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.0,1374.2,0,61,0,7.83,5011,0,Oakland,0,1,NA,37.80707,-122.29740100000001,1,20.0,1,4,None,21054,0,0,1,0,66,2,0.0,516.78,0.0,1374.2,0,0,94607
5972,0,1,0,0,15,1,1,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),55.0,757.1,1,73,21,17.19,3167,1,Emeryville,0,0,Cable,37.83726,-122.287648,0,57.2,0,0,Offer D,24589,1,1,0,0,15,1,159.0,257.85,0.0,757.1,0,0,94608
5973,1,0,0,0,64,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),104.4,6692.65,0,37,14,45.82,5617,0,Oakland,1,1,DSL,37.834340999999995,-122.26437,0,104.4,0,0,None,21097,0,0,0,1,64,1,93.7,2932.48,0.0,6692.65,0,1,94609
5974,1,0,1,1,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.05,218.5,0,55,0,13.83,2049,0,Oakland,0,1,NA,37.808731,-122.238708,1,20.05,3,7,None,29964,0,0,1,0,10,0,0.0,138.3,0.0,218.5,0,0,94610
5975,1,0,1,1,7,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.75,608.8,1,25,57,19.23,3807,1,Oakland,0,1,DSL,37.828416,-122.21600500000001,1,93.34,0,1,None,36517,1,1,1,0,7,5,347.0,134.61,26.02,608.8,1,0,94611
5976,1,0,0,0,29,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,34.3,1004.75,0,40,27,0.0,2555,0,Oakland,0,1,Fiber Optic,37.809014000000005,-122.26973899999999,0,34.3,0,0,None,11702,1,0,0,0,29,0,0.0,0.0,0.0,1004.75,0,1,94612
5977,1,0,0,0,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.65,1125.6,0,60,0,1.69,4193,0,Oakland,0,1,NA,37.84551,-122.23518100000001,0,20.65,0,0,None,15438,0,0,0,0,57,0,0.0,96.33,0.0,1125.6,0,0,94618
5978,0,0,0,0,46,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Mailed check,84.25,3847.6,0,37,21,43.27,3509,0,Oakland,0,0,Cable,37.787186,-122.14633,0,84.25,0,0,None,24518,0,0,0,0,46,0,80.8,1990.42,0.0,3847.6,0,1,94619
5979,1,0,0,0,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.65,978,0,62,0,23.17,5878,0,Oakland,0,1,NA,37.750553000000004,-122.197175,0,19.65,0,0,None,30751,0,0,0,0,53,0,0.0,1228.01,0.0,978.0,0,0,94621
5980,0,0,0,0,17,1,0,DSL,1,1,1,1,One year,0,Credit card (automatic),79.85,1387.35,0,45,22,12.69,5574,0,Berkeley,0,0,DSL,37.866009000000005,-122.28622800000001,0,79.85,0,0,None,15638,1,0,0,1,17,0,305.0,215.73,0.0,1387.35,0,0,94702
5981,0,0,1,1,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.2,746.05,0,54,0,26.84,2631,0,Berkeley,0,0,NA,37.863843,-122.27568400000001,1,20.2,1,9,None,19763,0,0,1,0,38,0,0.0,1019.92,0.0,746.05,0,0,94703
5982,1,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.8,304.6,0,49,0,5.54,5753,0,Berkeley,0,1,NA,37.871415999999996,-122.246597,0,19.8,0,0,None,21205,0,0,0,0,15,0,0.0,83.1,0.0,304.6,0,0,94704
5983,0,0,0,0,22,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,50.35,1098.85,0,51,22,0.0,2875,0,Berkeley,0,0,Cable,37.858897999999996,-122.24051200000001,0,50.35,0,0,None,12448,0,0,0,1,22,3,242.0,0.0,0.0,1098.85,0,0,94705
5984,1,0,1,0,14,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.15,1139.2,1,27,46,21.3,4550,1,Albany,0,1,Fiber Optic,37.890274,-122.29519199999999,1,88.55600000000003,0,1,None,15882,0,0,1,1,14,4,524.0,298.2,38.48,1139.2,1,0,94706
5985,0,0,1,0,57,1,1,DSL,0,1,1,0,One year,0,Bank transfer (automatic),74.6,4368.95,0,25,27,6.63,4546,0,Berkeley,1,0,Cable,37.897753,-122.27939099999999,1,74.6,0,2,None,11889,1,0,1,0,57,1,117.96,377.91,0.0,4368.95,1,1,94707
5986,1,1,0,0,11,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),79.15,827.7,0,80,15,26.84,3355,0,Berkeley,0,1,Fiber Optic,37.897743,-122.263124,0,79.15,0,0,Offer D,10737,0,0,0,1,11,4,0.0,295.24,0.0,827.7,0,1,94708
5987,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.35,20.35,0,62,0,30.09,4836,0,Berkeley,0,0,NA,37.878554,-122.26608999999999,1,20.35,3,9,None,10147,0,0,1,0,1,0,0.0,30.09,0.0,20.35,0,0,94709
5988,1,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),21.05,262.05,0,24,0,49.7,4843,0,Berkeley,0,1,NA,37.872902,-122.30370800000001,1,21.05,1,3,None,8157,0,0,1,0,12,0,0.0,596.4000000000002,0.0,262.05,1,0,94710
5989,1,1,1,0,3,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.6,279.55,1,70,30,32.31,3019,1,Richmond,0,1,DSL,37.945288,-122.383941,1,98.384,0,1,Offer E,28450,0,1,1,0,3,1,0.0,96.93,0.0,279.55,0,1,94801
5990,1,0,0,1,36,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,94.7,3512.5,0,55,18,21.3,4671,0,El Sobrante,0,1,Fiber Optic,37.963995000000004,-122.288296,0,94.7,1,0,None,25399,0,0,0,1,36,1,632.0,766.8000000000002,0.0,3512.5,0,0,94803
5991,1,0,0,0,16,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,94.25,1483.25,1,27,65,20.44,2827,1,Richmond,0,1,DSL,37.921034000000006,-122.341798,0,98.02,0,0,None,39089,0,1,0,1,16,2,964.0,327.04,0.0,1483.25,1,0,94804
5992,1,0,1,1,65,1,1,DSL,1,1,0,1,One year,0,Credit card (automatic),72.45,4653.85,1,24,56,26.75,4415,1,Richmond,1,1,DSL,37.941456,-122.320968,1,75.348,0,1,Offer B,13984,0,0,1,1,65,3,2606.0,1738.75,14.23,4653.85,1,0,94805
5993,1,0,0,0,2,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,74.95,151.75,0,54,16,3.76,3969,0,San Pablo,0,1,DSL,37.980269,-122.34263500000002,0,74.95,0,0,None,55720,0,0,0,0,2,0,0.0,7.52,0.0,151.75,0,1,94806
5994,0,0,0,0,42,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,105.2,4400.75,1,26,57,33.46,2317,1,San Rafael,1,0,Cable,37.972662,-122.491452,0,109.40799999999999,0,0,Offer B,40239,0,0,0,1,42,2,2508.0,1405.32,40.15,4400.75,1,0,94901
5995,1,0,1,1,72,1,0,Fiber optic,1,1,1,1,Two year,0,Bank transfer (automatic),111.95,8033.1,0,47,19,24.08,4004,0,San Rafael,1,1,Fiber Optic,38.018065,-122.546024,1,111.95,1,9,None,28403,1,0,1,1,72,1,1526.0,1733.7599999999998,0.0,8033.1,0,0,94903
5996,1,0,0,0,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.85,1253.65,0,29,0,14.17,4278,0,Greenbrae,0,1,NA,37.946616999999996,-122.563571,0,19.85,0,0,None,12010,0,0,0,0,62,1,0.0,878.54,0.0,1253.65,1,0,94904
5997,0,0,0,0,6,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.75,552.65,0,23,42,34.42,2370,0,Belvedere Tiburon,0,0,Fiber Optic,37.885628999999994,-122.46858,0,89.75,0,0,None,13065,0,0,0,0,6,1,232.0,206.52,0.0,552.65,1,0,94920
5998,1,0,1,0,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.05,1036,0,44,0,33.06,2964,0,Bodega,0,1,NA,38.343282,-122.9755,1,20.05,0,4,None,584,0,0,1,0,48,0,0.0,1586.88,0.0,1036.0,0,0,94922
5999,1,0,0,0,35,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,108.95,4025.5,0,42,23,20.07,5903,0,Bodega Bay,1,1,Cable,38.377165000000005,-123.037957,0,108.95,0,0,None,1785,1,0,0,1,35,0,0.0,702.45,0.0,4025.5,0,1,94923
6000,1,0,0,1,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.65,928.4,0,23,0,22.65,4279,0,Bolinas,0,1,NA,37.943087,-122.72379,0,19.65,2,0,None,1573,0,0,0,0,52,0,0.0,1177.8,0.0,928.4,1,0,94924
6001,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,24.9,24.9,0,37,13,0.0,5318,0,Corte Madera,0,0,Fiber Optic,37.924014,-122.51169399999999,0,24.9,0,0,None,9038,0,0,0,0,1,0,0.0,0.0,0.0,24.9,0,0,94925
6002,1,0,1,0,6,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,82.85,460.25,1,34,31,8.59,4458,1,Rohnert Park,0,1,Cable,38.347190000000005,-122.697822,1,86.164,0,3,None,42544,0,2,1,0,6,5,0.0,51.54,48.95,460.25,0,1,94928
6003,0,0,1,0,71,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),93.2,6506.15,0,38,23,12.12,4493,0,Dillon Beach,1,0,Fiber Optic,38.24458,-122.956268,1,93.2,0,8,None,330,1,1,1,1,71,1,0.0,860.52,0.0,6506.15,0,1,94929
6004,0,0,1,1,67,1,0,Fiber optic,1,1,0,0,One year,0,Bank transfer (automatic),84.8,5598.3,0,64,21,3.47,6072,0,Fairfax,1,0,Fiber Optic,37.971751,-122.611873,1,84.8,3,5,None,8486,0,0,1,0,67,0,0.0,232.49,0.0,5598.3,0,1,94930
6005,1,1,0,0,60,1,1,DSL,1,1,0,1,One year,1,Electronic check,71.75,4374.55,0,72,29,10.2,4964,0,Cotati,0,1,Cable,38.326215000000005,-122.71874199999999,0,71.75,0,0,None,7936,0,0,0,1,60,0,1269.0,612.0,0.0,4374.55,0,0,94931
6006,1,0,1,1,23,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),30.35,678.75,0,45,19,0.0,4960,0,Forest Knolls,0,1,Fiber Optic,38.010092,-122.68944199999999,1,30.35,1,2,Offer D,1025,1,0,1,0,23,0,129.0,0.0,0.0,678.75,0,0,94933
6007,1,0,0,1,39,0,No phone service,DSL,0,0,1,1,One year,0,Bank transfer (automatic),54.85,2191.7,0,31,29,0.0,3884,0,Inverness,1,1,DSL,38.099323,-122.945723,0,54.85,3,0,None,1004,1,0,0,1,39,3,0.0,0.0,0.0,2191.7,0,1,94937
6008,1,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.5,239.75,0,35,0,49.36,5471,0,Lagunitas,0,1,NA,38.021772,-122.691744,1,19.5,3,9,Offer D,821,0,0,1,0,15,0,0.0,740.4,0.0,239.75,0,0,94938
6009,1,1,1,0,53,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,103.85,5485.5,1,74,25,39.36,5860,1,Larkspur,1,1,DSL,37.937082000000004,-122.53236899999999,1,108.004,0,1,None,6773,0,1,1,0,53,2,1371.0,2086.08,0.0,5485.5,0,0,94939
6010,1,0,1,1,24,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.2,609.05,0,58,0,7.37,5865,0,Marshall,0,1,NA,38.129308,-122.83481499999999,1,24.2,3,1,None,406,0,1,1,0,24,2,0.0,176.88,0.0,609.05,0,0,94940
6011,0,0,1,1,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.35,683.75,0,20,0,2.68,2360,0,Mill Valley,0,0,NA,37.901371000000005,-122.572024,1,19.35,2,1,None,28727,0,0,1,0,37,2,0.0,99.16,0.0,683.75,1,0,94941
6012,0,0,1,1,5,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,83.6,404.2,1,54,25,7.0,4565,1,Novato,0,0,Fiber Optic,38.135897,-122.56368300000001,1,86.944,0,1,None,16429,0,0,1,1,5,1,101.0,35.0,24.44,404.2,0,0,94945
6013,0,1,1,0,50,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,100.65,5189.75,0,79,23,36.58,5791,0,Nicasio,0,0,Fiber Optic,38.065359,-122.665566,1,100.65,0,1,None,607,1,0,1,1,50,1,0.0,1829.0,0.0,5189.75,0,1,94946
6014,0,0,0,0,54,1,0,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),94.1,5060.9,0,23,42,48.97,4084,0,Novato,1,0,Fiber Optic,38.112165999999995,-122.63438400000001,0,94.1,0,0,None,24741,0,1,0,1,54,1,0.0,2644.38,0.0,5060.9,1,1,94947
6015,0,0,0,0,3,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,74.55,233.65,0,20,73,10.1,5125,0,Novato,0,0,Fiber Optic,38.067204,-122.524004,0,74.55,0,0,None,13361,0,1,0,0,3,1,171.0,30.3,0.0,233.65,1,0,94949
6016,1,0,0,0,68,1,1,Fiber optic,0,1,1,1,One year,0,Electronic check,108.45,7176.55,1,24,80,21.74,4454,1,Olema,1,1,Cable,38.052209000000005,-122.775567,0,112.788,0,0,Offer A,248,1,2,0,1,68,4,5741.0,1478.32,9.68,7176.55,1,0,94950
6017,1,0,0,0,5,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,56.15,291.45,0,23,71,26.86,5232,0,Penngrove,1,1,Fiber Optic,38.325599,-122.642352,0,56.15,0,0,None,3777,1,0,0,0,5,0,0.0,134.3,0.0,291.45,1,1,94951
6018,1,0,0,0,33,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.35,689.75,0,21,0,14.48,2507,0,Petaluma,0,1,NA,38.237018,-122.77871999999999,0,20.35,0,0,None,31930,0,0,0,0,33,0,0.0,477.84,0.0,689.75,1,0,94952
6019,0,0,0,0,41,1,1,DSL,0,1,1,1,One year,1,Electronic check,80.55,3263.9,0,51,12,6.16,4176,0,Petaluma,1,0,Fiber Optic,38.235021,-122.557332,0,80.55,0,0,None,35419,0,0,0,1,41,3,0.0,252.56,0.0,3263.9,0,1,94954
6020,0,0,1,1,34,0,No phone service,DSL,1,0,1,1,One year,0,Mailed check,61.25,1993.2,0,52,20,0.0,3607,0,Point Reyes Station,1,0,Fiber Optic,38.060264000000004,-122.830646,1,61.25,1,0,None,1885,1,0,0,1,34,1,399.0,0.0,0.0,1993.2,0,0,94956
6021,0,0,1,1,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.45,254.5,0,59,0,16.4,5417,0,San Anselmo,0,0,NA,37.99272,-122.575026,1,20.45,1,1,Offer D,16849,0,0,1,0,13,0,0.0,213.2,0.0,254.5,0,0,94960
6022,0,0,0,0,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),18.9,347.65,0,46,0,33.86,4277,0,San Geronimo,0,0,NA,38.004740000000005,-122.66371699999999,0,18.9,0,0,Offer D,548,0,0,0,0,20,3,0.0,677.2,0.0,347.65,0,0,94963
6023,0,1,0,0,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.6,967.9,0,66,0,47.46,4224,0,San Quentin,0,0,NA,37.942551,-122.491642,0,19.6,0,0,None,6448,0,0,0,0,51,1,0.0,2420.46,0.0,967.9,0,0,94964
6024,0,0,1,0,3,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),91.5,242.95,1,33,22,31.61,5646,1,Sausalito,0,0,Cable,37.848641,-122.51569199999999,1,95.16,0,1,None,11213,0,0,1,1,3,2,0.0,94.83,0.0,242.95,0,1,94965
6025,0,0,0,1,41,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),45.2,1841.9,0,58,28,38.94,4418,0,Stinson Beach,0,0,Cable,37.921137,-122.65756200000001,0,45.2,3,0,None,781,0,0,0,0,41,2,0.0,1596.54,0.0,1841.9,0,1,94970
6026,0,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.45,232.1,0,42,0,46.3,2783,0,Tomales,0,0,NA,38.240769,-122.90104099999999,0,19.45,0,0,Offer D,384,0,0,0,0,13,0,0.0,601.9,0.0,232.1,0,0,94971
6027,1,0,1,1,35,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.45,809.25,0,38,0,13.67,4873,0,Valley Ford,0,1,NA,38.339996,-122.935056,1,25.45,3,1,None,66,0,0,1,0,35,0,0.0,478.45,0.0,809.25,0,0,94972
6028,1,0,1,0,12,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Bank transfer (automatic),80.85,866.45,1,57,20,18.26,4306,1,Woodacre,0,1,DSL,38.005839,-122.638155,1,84.084,0,3,None,1449,1,0,1,0,12,4,173.0,219.12,23.72,866.45,0,0,94973
6029,1,0,0,0,4,1,0,Fiber optic,1,1,0,1,Month-to-month,1,Mailed check,94.9,360.55,0,25,41,11.5,3094,0,Alviso,0,1,Fiber Optic,37.449537,-121.994813,0,94.9,0,0,None,2147,1,0,0,1,4,1,148.0,46.0,0.0,360.55,1,0,95002
6030,0,0,0,0,43,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Bank transfer (automatic),49.05,2076.2,1,64,13,0.0,4044,1,Aptos,1,0,Cable,37.013471,-121.877877,0,51.012,0,0,Offer B,24227,0,0,0,1,43,2,270.0,0.0,20.29,2076.2,0,0,95003
6031,0,1,1,1,12,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,29.3,355.9,0,70,14,0.0,3353,0,Aromas,0,0,Fiber Optic,36.878364000000005,-121.62978100000001,1,29.3,1,1,Offer D,3373,1,0,1,0,12,1,50.0,0.0,0.0,355.9,0,0,95004
6032,1,1,1,0,68,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.3,7299.65,1,70,32,47.17,6284,1,Ben Lomond,1,1,Fiber Optic,37.078873,-122.09038600000001,1,109.512,0,1,None,6407,0,0,1,0,68,2,2336.0,3207.56,0.0,7299.65,0,0,95005
6033,1,1,0,0,25,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,88.95,2291.2,1,71,25,47.66,3878,1,Boulder Creek,0,1,Fiber Optic,37.171727000000004,-122.14296100000001,0,92.508,0,0,Offer C,10520,0,0,0,0,25,1,573.0,1191.5,0.0,2291.2,0,0,95006
6034,0,0,0,0,7,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.25,129.15,0,41,0,39.59,4208,0,Brookdale,0,0,NA,37.106902000000005,-122.10000600000001,0,20.25,0,0,None,1007,0,0,0,0,7,3,0.0,277.13,0.0,129.15,0,0,95007
6035,1,1,1,0,66,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,110.85,7491.75,1,66,14,48.87,4281,1,Campbell,1,1,DSL,37.279689000000005,-121.954567,1,115.284,0,1,None,44976,1,2,1,0,66,1,1049.0,3225.42,0.0,7491.75,0,0,95008
6036,0,0,1,0,53,1,0,Fiber optic,1,1,1,1,One year,0,Electronic check,110.5,5835.5,0,43,25,6.68,4135,0,Capitola,1,0,Fiber Optic,36.977025,-121.95286399999999,1,110.5,0,1,None,9673,1,0,1,1,53,1,145.89,354.04,0.0,5835.5,0,1,95010
6037,1,1,0,0,63,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),109.4,7031.45,0,68,20,26.11,5961,0,Castroville,1,1,Cable,36.784481,-121.759054,0,109.4,0,0,None,8582,0,0,0,1,63,0,1406.0,1644.93,0.0,7031.45,0,0,95012
6038,0,0,1,1,70,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.2,7723.9,1,21,53,16.78,5947,1,Cupertino,1,0,Cable,37.306612,-122.080621,1,118.76799999999999,0,1,Offer A,54431,1,0,1,1,70,3,0.0,1174.6,48.54,7723.9,1,1,95014
6039,1,1,1,0,27,0,No phone service,DSL,0,0,0,1,Month-to-month,0,Bank transfer (automatic),36.5,1032,1,68,28,0.0,4564,1,Davenport,0,1,DSL,37.114335,-122.23716200000001,1,37.96,0,1,Offer C,857,0,2,1,0,27,2,0.0,0.0,0.0,1032.0,0,1,95017
6040,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,70.75,70.75,1,56,9,26.0,3963,1,Felton,0,0,Cable,37.089110999999995,-122.06221299999999,0,73.58,0,0,None,8728,0,1,0,0,1,4,0.0,26.0,0.0,70.75,0,1,95018
6041,0,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,109.6,0,33,0,34.8,5252,0,Freedom,0,0,NA,36.936228,-121.785559,0,19.95,0,0,None,4753,0,0,0,0,5,0,0.0,174.0,0.0,109.6,0,0,95019
6042,0,1,1,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.6,727.8,0,77,0,25.35,5730,0,Gilroy,0,0,NA,37.03889,-121.52895500000001,1,19.6,0,1,None,49968,0,0,1,0,37,1,0.0,937.95,0.0,727.8,0,0,95020
6043,1,0,0,0,3,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Mailed check,40.15,130.75,1,19,29,0.0,4710,1,Escondido,1,1,DSL,33.141265000000004,-116.967221,0,41.756,0,0,None,48690,0,1,0,0,3,3,38.0,0.0,0.0,130.75,1,0,92027
6044,0,0,0,1,12,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.6,893,0,43,23,26.13,3280,0,Los Gatos,0,0,Cable,37.222842,-121.988727,0,76.6,1,0,Offer D,13290,0,0,0,0,12,2,205.0,313.56,0.0,893.0,0,0,95030
6045,0,0,1,1,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.6,763.1,0,60,0,36.72,4623,0,Los Gatos,0,0,NA,37.233034,-121.947427,1,19.6,2,1,None,24443,0,0,1,0,38,2,0.0,1395.36,0.0,763.1,0,0,95032
6046,0,0,0,0,9,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),85.3,781.4,0,64,8,48.38,5850,0,Los Gatos,1,0,Fiber Optic,37.160194,-121.94561100000001,0,85.3,0,0,None,10172,0,0,0,1,9,2,63.0,435.42,0.0,781.4,0,0,95033
6047,1,0,1,0,13,1,1,DSL,1,0,0,1,Month-to-month,1,Electronic check,65.85,902.25,0,56,4,14.32,2731,0,Milpitas,0,1,Fiber Optic,37.441931,-121.878502,1,65.85,0,1,Offer D,62848,0,0,1,1,13,3,3.61,186.16,0.0,902.25,0,1,95035
6048,1,1,1,0,29,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.45,2653.65,1,73,23,6.25,2233,1,Morgan Hill,0,1,Cable,37.161544,-121.649371,1,98.228,0,1,None,41707,0,6,1,0,29,1,610.0,181.25,0.0,2653.65,0,0,95037
6049,0,0,1,1,47,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.05,1016.7,0,52,0,1.44,3260,0,Moss Landing,0,0,NA,36.863303,-121.781632,1,20.05,1,1,None,899,0,0,1,0,47,0,0.0,67.67999999999999,0.0,1016.7,0,0,95039
6050,1,0,1,0,61,1,1,Fiber optic,1,0,1,0,Month-to-month,0,Bank transfer (automatic),99.4,5943.65,0,49,28,15.15,5404,0,Mount Hermon,1,1,Cable,37.051165999999995,-122.05619399999999,1,99.4,0,1,None,77,1,0,1,0,61,0,166.42,924.15,0.0,5943.65,0,1,95041
6051,1,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,275.7,0,22,0,4.13,3705,0,Paicines,0,1,NA,36.525703,-120.952122,0,20.0,0,0,Offer D,813,0,0,0,0,16,1,0.0,66.08,0.0,275.7,1,0,95043
6052,0,0,1,1,41,1,0,DSL,1,1,1,1,Two year,0,Electronic check,78.45,3126.45,0,20,69,32.29,5468,0,San Juan Bautista,0,0,DSL,36.810567999999996,-121.503022,1,78.45,2,1,None,3402,1,0,1,1,41,1,0.0,1323.89,0.0,3126.45,1,1,95045
6053,0,0,0,1,43,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Electronic check,25.1,1070.15,0,31,0,30.64,4797,0,San Martin,0,0,NA,37.084697,-121.606417,0,25.1,3,0,None,5671,0,0,0,0,43,2,0.0,1317.52,0.0,1070.15,0,0,95046
6054,0,0,1,1,36,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),97.35,3457.9,1,39,30,24.51,4544,1,Santa Clara,1,0,Fiber Optic,37.351214,-121.952417,1,101.244,0,3,None,36349,0,3,1,0,36,2,0.0,882.36,4.96,3457.9,0,1,95050
6055,0,0,0,0,6,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.0,340.4,0,27,58,37.57,2629,0,Santa Clara,0,0,Fiber Optic,37.348129,-121.98468999999999,0,55.0,0,0,None,52986,0,0,0,1,6,0,0.0,225.42,0.0,340.4,1,1,95051
6056,0,0,0,0,58,1,1,DSL,1,1,0,0,One year,1,Credit card (automatic),71.1,4299.2,0,56,7,42.33,5395,0,Santa Clara,1,0,Fiber Optic,37.393553999999995,-121.96511399999999,0,71.1,0,0,None,13031,1,0,0,0,58,0,301.0,2455.14,0.0,4299.2,0,0,95054
6057,1,0,0,0,19,1,0,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),61.55,1093.2,0,62,8,46.49,5831,0,Santa Cruz,0,1,Fiber Optic,36.993451,-122.098858,0,61.55,0,0,Offer D,43192,1,0,0,0,19,0,87.0,883.3100000000002,0.0,1093.2,0,0,95060
6058,1,0,1,0,11,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),45.9,521.9,0,54,6,12.95,3880,0,Santa Cruz,0,1,DSL,36.974575,-121.991149,1,45.9,0,1,Offer D,36631,0,0,1,0,11,0,3.13,142.45,0.0,521.9,0,1,95062
6059,0,0,0,0,39,0,No phone service,DSL,1,1,0,0,One year,1,Bank transfer (automatic),40.3,1630.4,0,37,19,0.0,3424,0,Santa Cruz,0,0,Fiber Optic,37.007882,-122.065975,0,40.3,0,0,None,4563,1,0,0,0,39,0,310.0,0.0,0.0,1630.4,0,0,95064
6060,0,1,0,0,8,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,87.1,713.6,0,80,28,39.01,3950,0,Santa Cruz,0,0,Fiber Optic,37.031403999999995,-121.98186499999998,0,87.1,0,0,None,8365,0,0,0,0,8,0,200.0,312.08,0.0,713.6,0,0,95065
6061,0,0,0,1,26,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,49.5,1265.65,0,53,19,16.34,4196,0,Scotts Valley,0,0,DSL,37.070177,-122.010077,0,49.5,1,0,None,14574,0,0,0,0,26,2,24.05,424.84,0.0,1265.65,0,1,95066
6062,0,1,0,0,53,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),73.8,4003.85,0,75,15,16.74,6469,0,Saratoga,0,0,Cable,37.257771999999996,-122.051824,0,73.8,0,0,None,30589,0,0,0,0,53,0,60.06,887.2199999999998,0.0,4003.85,0,1,95070
6063,0,0,1,1,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.2,1401.4,0,38,0,38.63,5261,0,Soquel,0,0,NA,37.023669,-121.94646100000001,1,19.2,3,1,None,9823,0,1,1,0,70,2,0.0,2704.100000000001,0.0,1401.4,0,0,95073
6064,1,0,0,0,1,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Mailed check,45.3,45.3,1,34,20,0.0,4954,1,Watsonville,0,1,DSL,36.931653999999995,-121.75238300000001,0,47.111999999999995,0,0,None,81141,0,1,0,1,1,4,0.0,0.0,0.0,45.3,0,0,95076
6065,1,0,0,0,59,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.0,1510.5,0,25,0,25.89,5537,0,San Jose,0,1,NA,37.34667,-121.91001899999999,0,25.0,0,0,None,18197,0,0,0,0,59,1,0.0,1527.51,0.0,1510.5,1,0,95110
6066,1,0,0,0,2,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,94.95,178.1,1,61,2,26.05,4493,1,San Jose,1,1,DSL,37.284265000000005,-121.827673,0,98.74799999999999,0,0,None,57748,0,1,0,1,2,1,4.0,52.1,0.0,178.1,0,0,95111
6067,1,0,0,0,7,0,No phone service,DSL,1,0,0,0,One year,0,Mailed check,35.3,264.8,0,47,14,0.0,3463,0,San Jose,1,1,DSL,37.343827000000005,-121.883119,0,35.3,0,0,None,52334,0,0,0,0,7,3,0.0,0.0,0.0,264.8,0,1,95112
6068,0,0,0,1,12,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.55,480.6,1,33,18,5.16,4162,1,San Jose,0,0,DSL,37.333851,-121.891147,0,46.332,1,0,None,561,0,1,0,0,12,4,87.0,61.92,18.21,480.6,0,0,95113
6069,1,0,1,1,59,1,0,DSL,0,1,1,1,One year,0,Credit card (automatic),76.75,4541.9,0,63,19,15.94,5918,0,San Jose,1,1,Fiber Optic,37.350284,-121.852855,1,76.75,2,1,None,51706,1,0,1,1,59,2,0.0,940.46,0.0,4541.9,0,1,95116
6070,1,0,1,1,61,1,1,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),81.0,4976.15,0,27,41,32.96,4151,0,San Jose,1,1,Fiber Optic,37.311088,-121.961786,1,81.0,3,1,None,29914,1,0,1,1,61,0,2040.0,2010.56,0.0,4976.15,1,0,95117
6071,1,0,1,1,72,1,1,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),105.55,7542.25,0,22,59,8.33,4331,0,San Jose,1,1,DSL,37.255479,-121.88983799999998,1,105.55,3,4,None,31926,0,0,1,1,72,1,0.0,599.76,0.0,7542.25,1,1,95118
6072,0,0,1,1,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,18.8,251.25,0,27,0,16.74,2333,0,San Jose,0,0,NA,37.233226,-121.78809,1,18.8,1,6,Offer D,10155,0,0,1,0,13,1,0.0,217.62,0.0,251.25,1,0,95119
6073,0,0,1,1,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,24.9,1595.5,0,50,0,19.23,5038,0,San Jose,0,0,NA,37.186141,-121.843554,1,24.9,1,6,None,37090,0,0,1,0,64,0,0.0,1230.72,0.0,1595.5,0,0,95120
6074,1,0,1,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,23.45,23.45,1,55,23,0.0,4517,1,San Jose,0,1,DSL,37.304681,-121.809955,1,24.388,0,3,Offer E,37127,0,0,1,0,1,3,0.0,0.0,0.0,23.45,0,0,95121
6075,0,0,0,0,10,1,0,DSL,0,1,0,1,One year,0,Mailed check,64.9,685.55,0,54,5,37.45,4883,0,San Jose,0,0,Cable,37.32886,-121.83456699999999,0,64.9,0,0,Offer D,59841,1,0,0,1,10,0,3.43,374.5,0.0,685.55,0,1,95122
6076,0,0,1,1,65,1,0,DSL,1,1,0,0,One year,0,Bank transfer (automatic),61.35,3874.1,0,55,19,19.25,6354,0,San Jose,1,0,Fiber Optic,37.238758000000004,-121.828375,1,61.35,2,0,Offer B,59632,0,0,0,0,65,1,0.0,1251.25,0.0,3874.1,0,1,95123
6077,0,0,1,0,62,1,1,Fiber optic,1,1,1,1,Two year,0,Mailed check,113.95,6891.4,0,21,51,42.68,6193,0,San Jose,1,0,DSL,37.257063,-121.92303700000001,1,113.95,0,3,Offer B,45257,1,0,1,1,62,0,0.0,2646.16,0.0,6891.4,1,1,95124
6078,0,0,1,0,55,1,1,DSL,1,1,1,1,One year,1,Electronic check,90.15,4916.95,0,20,53,47.46,4712,0,San Jose,1,0,DSL,37.294926000000004,-121.89476299999998,1,90.15,0,8,Offer B,46185,1,0,1,1,55,0,0.0,2610.3,0.0,4916.95,1,1,95125
6079,0,0,1,0,25,1,1,DSL,0,1,0,0,Month-to-month,0,Electronic check,54.1,1373,0,29,59,12.12,5701,0,San Jose,0,0,Cable,37.327069,-121.91681899999999,1,54.1,0,8,None,27023,0,1,1,0,25,1,0.0,303.0,0.0,1373.0,1,1,95126
6080,1,0,0,0,1,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Mailed check,29.7,29.7,1,30,76,0.0,3383,1,San Jose,0,1,Cable,37.375156,-121.79586699999999,0,30.888,0,0,Offer E,60620,0,4,0,0,1,4,0.0,0.0,0.0,29.7,0,1,95127
6081,1,0,0,0,1,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),49.8,49.8,0,55,13,38.21,2978,0,San Jose,0,1,Fiber Optic,37.316146,-121.93628500000001,0,49.8,0,0,None,32804,0,0,0,0,1,1,0.0,38.21,0.0,49.8,0,1,95128
6082,0,0,1,0,59,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,101.1,6039.9,1,21,53,9.23,4160,1,San Jose,0,0,Cable,37.305622,-122.000887,1,105.144,0,4,Offer B,37570,0,1,1,1,59,4,3201.0,544.57,0.0,6039.9,1,0,95129
6083,1,1,1,1,64,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.4,1548.65,0,69,0,37.09,4772,0,San Jose,0,1,NA,37.277592,-121.98647700000001,1,24.4,1,9,None,13481,0,0,1,0,64,0,0.0,2373.76,0.0,1548.65,0,0,95130
6084,1,0,1,0,36,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.0,3440.25,0,50,6,5.99,3057,0,San Jose,0,1,Cable,37.387027,-121.897775,1,95.0,0,3,None,26389,0,0,1,1,36,1,206.0,215.64,0.0,3440.25,0,0,95131
6085,0,0,0,0,3,1,1,DSL,0,0,0,0,Month-to-month,1,Mailed check,50.65,151.3,1,51,3,22.56,2876,1,San Jose,0,0,Fiber Optic,37.424655,-121.74841,0,52.676,0,0,Offer E,40568,0,0,0,0,3,5,0.0,67.67999999999999,0.0,151.3,0,1,95132
6086,1,0,1,0,61,1,1,DSL,1,0,0,1,Two year,1,Mailed check,69.9,4226.7,0,37,4,4.69,5117,0,San Jose,1,1,Fiber Optic,37.371862,-121.860349,1,69.9,0,1,Offer B,26032,0,0,1,1,61,0,169.0,286.0900000000001,0.0,4226.7,0,0,95133
6087,1,0,0,1,26,0,No phone service,DSL,0,1,1,0,One year,1,Bank transfer (automatic),39.95,1023.75,0,32,58,0.0,2715,0,San Jose,0,1,Cable,37.42765,-121.945416,0,39.95,3,0,None,9657,0,0,0,0,26,2,594.0,0.0,0.0,1023.75,0,0,95134
6088,0,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.4,55.4,1,37,4,13.01,2294,1,San Jose,0,0,DSL,37.28682,-121.723877,0,57.61600000000001,0,0,Offer E,15798,0,2,0,1,1,1,0.0,13.01,0.0,55.4,0,0,95135
6089,0,1,1,0,1,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,90.6,90.6,1,77,33,13.02,2905,1,San Jose,0,0,DSL,37.270938,-121.851046,1,94.22399999999999,0,1,Offer E,36944,0,1,1,0,1,2,0.0,13.02,0.0,90.6,0,1,95136
6090,1,0,1,1,68,1,0,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),103.25,7074.4,0,51,29,21.86,4751,0,San Jose,1,1,Cable,37.246064000000004,-121.749494,1,103.25,2,2,None,14792,0,0,1,1,68,0,0.0,1486.48,0.0,7074.4,0,1,95138
6091,1,1,1,0,2,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,86.85,156.35,1,73,12,4.19,5204,1,San Jose,0,1,DSL,37.218705,-121.762429,1,90.324,0,3,None,7023,0,3,1,0,2,2,19.0,8.38,0.0,156.35,0,0,95139
6092,0,0,1,0,72,1,1,Fiber optic,1,1,0,0,Two year,1,Bank transfer (automatic),94.25,6849.75,0,39,17,11.02,6295,0,Mount Hamilton,1,0,Cable,37.382909000000005,-121.634151,1,94.25,0,8,None,38,1,0,1,0,72,1,1164.0,793.4399999999998,0.0,6849.75,0,0,95140
6093,0,0,1,0,71,0,No phone service,DSL,0,0,0,1,Two year,1,Electronic check,47.05,3263.6,0,59,6,0.0,6302,0,San Jose,1,0,Cable,37.339533,-121.777179,1,47.05,0,4,None,44103,1,0,1,1,71,2,196.0,0.0,0.0,3263.6,0,0,95148
6094,1,0,0,0,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.55,1252.85,0,56,0,12.99,4565,0,Stockton,0,1,NA,37.959706,-121.287669,0,20.55,0,0,Offer B,7071,0,1,0,0,57,3,0.0,740.4300000000002,0.0,1252.85,0,0,95202
6095,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.65,67.55,0,20,0,18.28,4925,0,Stockton,0,1,NA,37.954089,-121.329761,0,19.65,0,0,Offer E,16357,0,0,0,0,4,1,0.0,73.12,0.0,67.55,1,0,95203
6096,0,1,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.2,70.2,0,69,12,22.34,2422,0,Stockton,0,0,Fiber Optic,37.974498,-121.31956799999999,0,70.2,0,0,None,30476,0,1,0,0,1,2,0.0,22.34,0.0,70.2,0,1,95204
6097,1,0,1,1,72,1,1,DSL,1,1,0,1,Two year,0,Credit card (automatic),81.0,5750,0,22,59,2.73,4237,0,Stockton,1,1,DSL,37.965695000000004,-121.260051,1,81.0,3,8,None,34138,1,0,1,1,72,0,0.0,196.56,0.0,5750.0,1,1,95205
6098,1,0,1,1,21,1,1,DSL,1,0,1,1,One year,1,Bank transfer (automatic),75.9,1549.75,0,42,23,31.55,3503,0,Stockton,0,1,Fiber Optic,37.902421999999994,-121.44002900000001,1,75.9,3,6,None,49657,0,0,1,1,21,2,35.64,662.5500000000002,0.0,1549.75,0,1,95206
6099,0,0,1,1,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.7,1810.55,0,42,0,19.49,5187,0,Stockton,0,0,NA,38.002125,-121.324979,1,24.7,1,1,None,49965,0,0,1,0,71,0,0.0,1383.79,0.0,1810.55,0,0,95207
6100,0,1,1,0,29,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),99.05,2952.85,1,65,7,22.33,3179,1,Stockton,1,0,DSL,38.044523,-121.34804799999999,1,103.012,0,1,None,30814,0,0,1,1,29,0,207.0,647.5699999999998,0.0,2952.85,0,0,95209
6101,0,1,0,0,69,1,1,Fiber optic,1,0,1,1,Two year,0,Credit card (automatic),110.25,7467.55,0,72,27,23.4,4948,0,Stockton,1,0,Fiber Optic,38.033219,-121.29743300000001,0,110.25,0,0,None,40611,1,0,0,1,69,0,201.62,1614.6,0.0,7467.55,0,1,95210
6102,0,0,1,0,64,1,1,DSL,1,0,1,1,Two year,1,Credit card (automatic),85.0,5484.4,0,41,2,11.85,5472,0,Stockton,1,0,DSL,38.049457000000004,-121.21653,1,85.0,0,5,Offer B,6951,1,1,1,1,64,2,110.0,758.4,0.0,5484.4,0,0,95212
6103,1,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.75,294.9,0,48,0,24.79,5433,0,Stockton,0,1,NA,37.946282000000004,-121.139499,0,19.75,0,0,None,23789,0,0,0,0,16,0,0.0,396.64,0.0,294.9,0,0,95215
6104,0,0,0,0,4,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,23.9,97.5,0,33,0,6.36,5685,0,Stockton,0,0,NA,38.029728999999996,-121.387999,0,23.9,0,0,Offer E,19109,0,0,0,0,4,0,0.0,25.44,0.0,97.5,0,0,95219
6105,0,0,0,0,52,1,1,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),111.25,5916.45,1,20,57,33.69,4861,1,Acampo,0,0,Cable,38.200231,-121.23503400000001,0,115.7,0,0,Offer B,6317,1,0,0,1,52,1,3372.0,1751.88,1.27,5916.45,1,0,95220
6106,1,0,0,0,2,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,55.1,113.35,1,19,57,5.33,4235,1,Angels Camp,1,1,DSL,38.071327000000004,-120.632221,0,57.303999999999995,0,0,Offer E,4264,0,0,0,0,2,4,65.0,10.66,0.0,113.35,1,0,95222
6107,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,19.95,0,44,0,27.08,5916,0,Arnold,0,1,NA,38.321529999999996,-120.23635800000001,0,19.95,0,0,Offer E,5159,0,0,0,0,1,0,0.0,27.08,0.0,19.95,0,0,95223
6108,1,0,0,0,18,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,25.15,476.8,0,32,8,0.0,2675,0,Avery,0,1,Fiber Optic,38.208335999999996,-120.33993799999999,0,25.15,0,0,None,115,0,0,0,0,18,2,0.0,0.0,0.0,476.8,0,1,95224
6109,0,0,0,0,2,1,1,DSL,0,1,0,0,Month-to-month,0,Mailed check,54.15,101.65,0,47,7,21.3,3527,0,Burson,0,0,DSL,38.183918,-120.898817,0,54.15,0,0,Offer E,27,0,0,0,0,2,2,0.0,42.6,0.0,101.65,0,1,95225
6110,0,0,1,0,19,1,0,DSL,0,1,0,1,Month-to-month,1,Mailed check,59.8,1130.85,0,20,48,8.3,3652,0,Campo Seco,0,0,Fiber Optic,38.233878999999995,-120.86166599999999,1,59.8,0,3,None,75,0,1,1,1,19,1,0.0,157.70000000000005,0.0,1130.85,1,1,95226
6111,0,0,0,0,40,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Bank transfer (automatic),83.85,3532.25,0,50,20,33.66,4294,0,Clements,0,0,DSL,38.227284999999995,-121.02788999999999,0,83.85,0,0,Offer B,722,0,0,0,1,40,2,706.0,1346.4,0.0,3532.25,0,0,95227
6112,0,1,1,1,66,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,104.9,6891.45,0,67,30,39.38,4892,0,Copperopolis,1,0,DSL,37.943954,-120.67108,1,104.9,1,6,None,2633,0,0,1,1,66,1,2067.0,2599.080000000001,0.0,6891.45,0,0,95228
6113,1,0,0,0,21,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,75.3,1570.7,0,25,51,3.26,2847,0,Farmington,0,1,Fiber Optic,37.956963,-120.863055,0,75.3,0,0,None,596,0,0,0,0,21,1,80.11,68.46,0.0,1570.7,1,1,95230
6114,1,0,0,0,8,1,0,DSL,0,1,1,0,Month-to-month,1,Electronic check,66.65,520.95,0,41,27,30.8,3804,0,French Camp,0,1,Fiber Optic,37.873283,-121.29203400000002,0,66.65,0,0,Offer E,5094,1,0,0,0,8,0,0.0,246.4,0.0,520.95,0,1,95231
6115,0,0,1,1,72,1,0,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),109.5,7854.9,0,38,19,32.23,6419,0,Glencoe,1,0,Fiber Optic,38.358464,-120.57930400000001,1,109.5,1,3,None,21,1,0,1,1,72,0,149.24,2320.56,0.0,7854.9,0,1,95232
6116,0,0,0,0,48,1,1,DSL,0,1,1,0,One year,1,Bank transfer (automatic),73.85,3581.4,0,49,3,21.39,4740,0,Hathaway Pines,1,0,Cable,38.184914,-120.364085,0,73.85,0,0,Offer B,335,1,0,0,0,48,2,0.0,1026.72,0.0,3581.4,0,1,95233
6117,1,0,0,0,69,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.3,1447.9,0,54,0,17.74,5028,0,Linden,0,1,NA,38.047746000000004,-121.030499,0,19.3,0,0,None,3148,0,0,0,0,69,1,0.0,1224.06,0.0,1447.9,0,0,95236
6118,1,0,0,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,118.2,8547.15,0,60,27,36.49,4886,0,Lockeford,1,1,Fiber Optic,38.166790999999996,-121.14206999999999,0,118.2,0,0,None,3205,1,0,0,1,72,0,2308.0,2627.28,0.0,8547.15,0,0,95237
6119,0,0,0,0,14,1,0,DSL,0,1,0,0,One year,0,Credit card (automatic),51.45,727.85,0,64,12,24.04,4298,0,Lodi,0,0,DSL,38.123544,-121.15907800000001,0,51.45,0,0,None,45755,0,1,0,0,14,2,87.0,336.56,0.0,727.85,0,0,95240
6120,1,0,0,0,6,1,0,DSL,0,1,1,0,Month-to-month,0,Electronic check,59.45,357.6,0,58,8,10.88,2393,0,Lodi,0,1,DSL,38.128087,-121.4078,0,59.45,0,0,None,22073,0,0,0,0,6,1,29.0,65.28,0.0,357.6,0,0,95242
6121,0,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.5,159.35,0,48,0,17.2,5206,0,Mokelumne Hill,0,0,NA,38.304194,-120.592431,1,19.5,3,6,None,2718,0,1,1,0,8,3,0.0,137.6,0.0,159.35,0,0,95245
6122,0,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.55,280.85,0,21,0,42.42,4947,0,Mountain Ranch,0,0,NA,38.264262,-120.515133,0,19.55,0,0,None,1692,0,0,0,0,17,0,0.0,721.14,0.0,280.85,1,0,95246
6123,1,0,0,0,65,1,1,Fiber optic,1,0,0,1,One year,0,Electronic check,93.55,6069.25,0,50,16,2.72,5774,0,Murphys,0,1,DSL,38.147852,-120.440124,0,93.55,0,0,Offer B,4353,1,0,0,1,65,1,0.0,176.8,0.0,6069.25,0,1,95247
6124,0,0,1,1,57,1,0,DSL,1,0,0,0,One year,1,Mailed check,59.3,3274.35,0,54,24,18.85,6287,0,San Andreas,1,0,Fiber Optic,38.196496999999994,-120.61688999999998,1,59.3,1,6,Offer B,3930,1,0,1,0,57,1,0.0,1074.45,0.0,3274.35,0,1,95249
6125,1,0,1,0,13,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),102.25,1359,1,36,31,30.55,2003,1,Sheep Ranch,1,1,Cable,38.244806,-120.417301,1,106.34,0,1,None,88,0,0,1,1,13,0,421.0,397.15,0.0,1359.0,0,0,95250
6126,1,1,0,0,19,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),95.9,1777.9,1,65,4,32.77,2851,1,Vallecito,1,1,Fiber Optic,38.055562,-120.456298,0,99.736,0,0,Offer D,460,0,0,0,1,19,0,71.0,622.6300000000001,0.0,1777.9,0,0,95251
6127,0,0,1,0,56,1,1,Fiber optic,1,1,1,1,One year,0,Bank transfer (automatic),109.8,6109.65,0,54,21,37.76,5648,0,Valley Springs,1,0,DSL,38.156971,-120.849231,1,109.8,0,9,Offer B,11266,0,0,1,1,56,3,0.0,2114.56,0.0,6109.65,0,1,95252
6128,0,0,1,0,14,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,78.1,1122.4,0,50,16,4.45,3157,0,Wallace,0,0,Fiber Optic,38.192608,-120.957842,1,78.1,0,7,None,304,0,0,1,1,14,1,0.0,62.3,0.0,1122.4,0,1,95254
6129,1,0,1,0,52,0,No phone service,DSL,1,0,0,1,Month-to-month,1,Electronic check,39.9,2020.9,0,47,26,0.0,6371,0,West Point,0,1,Fiber Optic,38.41935,-120.469545,1,39.9,0,1,None,2198,0,0,1,1,52,2,0.0,0.0,0.0,2020.9,0,1,95255
6130,0,0,0,0,58,1,0,DSL,1,1,0,0,Two year,1,Credit card (automatic),64.9,3795.45,0,56,16,29.47,5040,0,Wilseyville,1,0,Cable,38.392686,-120.415951,0,64.9,0,0,None,435,1,0,0,0,58,0,607.0,1709.26,0.0,3795.45,0,0,95257
6131,0,1,0,0,47,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,95.05,4504.55,1,78,12,14.22,5214,1,Woodbridge,0,0,Fiber Optic,38.169605,-121.31096399999998,0,98.852,0,0,None,4176,1,0,0,0,47,1,541.0,668.34,0.0,4504.55,0,0,95258
6132,0,0,0,0,67,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),53.4,3579.15,0,61,11,0.0,5990,0,Atwater,1,0,DSL,37.321233,-120.65635400000001,0,53.4,0,0,None,27808,1,0,0,1,67,2,0.0,0.0,0.0,3579.15,0,1,95301
6133,1,0,0,0,2,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),24.9,49.7,0,22,48,0.0,4033,0,Ballico,0,1,DSL,37.4695,-120.672724,0,24.9,0,0,None,809,0,0,0,0,2,0,0.0,0.0,0.0,49.7,1,1,95303
6134,1,1,0,0,6,1,0,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),44.7,276.5,0,69,7,19.74,4270,0,Big Oak Flat,0,1,Cable,37.818589,-120.25699499999999,0,44.7,0,0,Offer E,167,0,0,0,0,6,0,0.0,118.44,0.0,276.5,0,1,95305
6135,1,0,1,1,71,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),114.0,8175.9,0,25,59,25.45,5600,0,Catheys Valley,1,1,Fiber Optic,37.394411,-120.12726200000002,1,114.0,1,0,None,986,1,0,0,1,71,1,0.0,1806.95,0.0,8175.9,1,1,95306
6136,0,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.25,890.35,0,42,0,27.65,3879,0,Ceres,0,0,NA,37.553469,-120.952825,1,20.25,1,7,None,32881,0,0,1,0,46,1,0.0,1271.9,0.0,890.35,0,0,95307
6137,0,0,0,0,5,1,0,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),53.85,259.8,1,34,24,24.32,5435,1,Columbia,0,0,Fiber Optic,38.085839,-120.37855,0,56.00400000000001,0,0,Offer E,2144,1,1,0,0,5,1,0.0,121.6,22.96,259.8,0,1,95310
6138,1,1,1,0,67,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Bank transfer (automatic),83.85,5588.8,0,66,20,44.9,5261,0,Coulterville,0,1,Cable,37.722127,-120.110174,1,83.85,0,10,None,2271,0,0,1,0,67,0,111.78,3008.3,0.0,5588.8,0,1,95311
6139,1,0,0,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.2,50.6,0,36,0,18.43,3594,0,Cressey,0,1,NA,37.420273,-120.66526999999999,0,20.2,3,0,None,55,0,0,0,0,3,1,0.0,55.29,0.0,50.6,0,0,95312
6140,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.95,58,0,60,0,2.69,5949,0,Crows Landing,0,0,NA,37.435664,-121.04905600000001,0,19.95,0,0,None,1508,0,0,0,0,3,2,0.0,8.07,0.0,58.0,0,0,95313
6141,1,1,1,0,52,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,104.2,5568.35,1,69,25,37.6,5648,1,Delhi,1,1,Fiber Optic,37.422961,-120.76549299999999,1,108.368,0,0,None,10159,0,0,0,1,52,1,1392.0,1955.2,0.0,5568.35,0,0,95315
6142,0,0,1,0,42,1,1,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.25,2203.65,1,30,45,10.79,4873,1,Denair,0,0,DSL,37.524721,-120.757977,1,52.26000000000001,0,2,Offer B,5513,0,1,1,0,42,2,992.0,453.18,28.49,2203.65,0,0,95316
6143,1,0,1,1,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,20.35,938.95,0,40,0,26.98,6391,0,El Nido,0,1,NA,37.127386,-120.506422,1,20.35,2,9,None,808,0,0,1,0,50,0,0.0,1349.0,0.0,938.95,0,0,95317
6144,1,1,1,0,23,1,0,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,90.0,2024.1,0,70,20,31.53,4999,0,El Portal,0,1,Fiber Optic,37.654551,-119.822984,1,90.0,0,3,Offer D,579,0,0,1,0,23,1,0.0,725.19,0.0,2024.1,0,1,95318
6145,0,0,1,1,67,0,No phone service,DSL,1,1,1,0,Two year,0,Credit card (automatic),54.2,3623.95,0,29,51,0.0,5261,0,Escalon,1,0,DSL,37.818543,-121.00690700000001,1,54.2,2,2,None,11474,1,1,1,0,67,2,0.0,0.0,0.0,3623.95,1,1,95320
6146,0,0,0,0,25,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,99.5,2369.05,1,35,9,48.42,5932,1,Groveland,1,0,Cable,37.902968,-119.66754399999999,0,103.48,0,0,None,3680,0,2,0,1,25,1,213.0,1210.5,19.5,2369.05,0,0,95321
6147,0,1,1,0,39,1,0,Fiber optic,1,1,1,1,One year,0,Mailed check,99.1,3877.95,0,77,18,9.13,4599,0,Gustine,0,0,Fiber Optic,37.147197999999996,-121.12016100000001,1,99.1,0,6,None,7872,0,0,1,0,39,0,69.8,356.07000000000005,0.0,3877.95,0,1,95322
6148,0,0,0,0,69,1,1,DSL,1,1,0,0,Two year,1,Mailed check,66.9,4577.9,0,46,7,13.91,5059,0,Hickman,0,0,Fiber Optic,37.605926000000004,-120.69955,0,66.9,0,0,Offer A,1055,1,0,0,0,69,2,32.05,959.79,0.0,4577.9,0,1,95323
6149,0,0,0,0,1,0,No phone service,DSL,0,0,0,0,One year,0,Mailed check,25.85,25.85,0,50,18,0.0,4467,0,Hilmar,0,0,DSL,37.394535999999995,-120.89074699999999,0,25.85,0,0,None,7177,0,0,0,0,1,0,0.0,0.0,0.0,25.85,0,1,95324
6150,1,0,0,0,32,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,91.05,2871.5,0,40,24,47.3,2716,0,Hornitos,0,1,DSL,37.479926,-120.230424,0,91.05,0,0,None,128,0,0,0,1,32,0,0.0,1513.6,0.0,2871.5,0,1,95325
6151,0,0,0,0,9,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,71.0,672.55,1,49,10,24.52,2236,1,Hughson,0,0,Cable,37.5923,-120.85328799999999,0,73.84,0,0,None,6822,0,1,0,0,9,1,67.0,220.68,8.35,672.55,0,0,95326
6152,0,0,0,0,16,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),93.2,1573.7,1,40,8,40.76,5497,1,Jamestown,1,0,DSL,37.84771,-120.486589,0,96.928,0,0,None,9559,0,0,0,1,16,0,126.0,652.16,35.7,1573.7,0,0,95327
6153,1,0,1,1,60,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.95,1270.55,0,45,0,32.12,4425,0,Keyes,0,1,NA,37.555631,-120.911653,1,20.95,2,9,None,2130,0,0,1,0,60,0,0.0,1927.2,0.0,1270.55,0,0,95328
6154,0,0,1,1,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),109.2,7711.45,0,40,14,44.03,6130,0,La Grange,1,0,Fiber Optic,37.666587,-120.41151699999999,1,109.2,1,4,Offer A,1749,1,0,1,1,72,0,1080.0,3170.16,0.0,7711.45,0,0,95329
6155,1,0,1,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.35,126.05,1,53,0,31.76,3864,1,Lathrop,0,1,NA,37.808209999999995,-121.308401,1,19.35,0,0,Offer E,10834,0,0,0,0,5,1,0.0,158.8,0.0,126.05,0,0,95330
6156,0,1,0,0,26,1,0,Fiber optic,1,0,1,0,Month-to-month,1,Credit card (automatic),85.8,2193.65,0,71,7,33.74,5700,0,Le Grand,0,0,Fiber Optic,37.249377,-120.249581,0,85.8,0,0,None,3256,0,0,0,0,26,2,154.0,877.24,0.0,2193.65,0,0,95333
6157,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.85,64.55,1,29,0,32.01,2158,1,Livingston,0,1,NA,37.361987,-120.74839399999999,0,19.85,0,0,Offer E,12672,0,0,0,0,3,1,0.0,96.03,0.0,64.55,1,0,95334
6158,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.65,31.2,0,55,0,7.8,4841,0,Long Barn,0,1,NA,38.109125,-120.078597,0,19.65,0,0,None,683,0,0,0,0,2,1,0.0,15.6,0.0,31.2,0,0,95335
6159,0,0,0,1,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.5,38.25,0,44,0,31.01,4486,0,Manteca,0,0,NA,37.830267,-121.20101799999999,0,20.5,3,0,None,36738,0,0,0,0,2,0,0.0,62.02,0.0,38.25,0,0,95336
6160,0,0,0,0,36,1,1,DSL,1,0,1,1,One year,1,Credit card (automatic),89.65,3348.1,0,29,59,44.7,4844,0,Manteca,1,0,DSL,37.750822,-121.238423,0,89.65,0,0,None,19867,1,0,0,1,36,0,1975.0,1609.2,0.0,3348.1,1,0,95337
6161,1,0,0,0,7,1,0,Fiber optic,1,0,0,0,Month-to-month,0,Mailed check,74.35,533.6,0,48,23,1.67,2463,0,Mariposa,0,1,Cable,37.526790999999996,-119.99436999999999,0,74.35,0,0,None,10226,0,0,0,0,7,1,0.0,11.69,0.0,533.6,0,1,95338
6162,0,1,1,0,60,0,No phone service,DSL,0,1,1,1,Two year,1,Credit card (automatic),49.45,2907.55,0,70,22,0.0,4277,0,Merced,0,0,DSL,37.255637,-120.49353700000002,1,49.45,0,3,None,59289,0,0,1,0,60,1,0.0,0.0,0.0,2907.55,0,1,95340
6163,0,0,1,0,19,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,89.1,1620.8,0,30,52,45.37,3624,0,Midpines,0,0,DSL,37.581496,-119.97276200000002,1,89.1,0,1,None,433,0,0,1,1,19,0,0.0,862.03,0.0,1620.8,0,1,95345
6164,1,1,1,0,45,1,1,DSL,1,0,0,1,Two year,0,Credit card (automatic),75.15,3480.35,0,77,22,9.39,5837,0,Mi Wuk Village,1,1,Cable,38.121601,-120.13391499999999,1,75.15,0,4,None,1278,1,0,1,0,45,1,766.0,422.55,0.0,3480.35,0,0,95346
6165,1,1,0,0,4,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.65,293.85,0,69,12,6.18,4510,0,Merced,0,1,Fiber Optic,37.40122,-120.514191,0,70.65,0,0,Offer E,23100,0,0,0,0,4,0,35.0,24.72,0.0,293.85,0,0,95348
6166,0,0,1,1,31,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,104.2,3243.45,1,51,14,3.73,5000,1,Modesto,1,0,DSL,37.671806,-121.007575,1,108.368,0,4,None,52872,1,2,1,1,31,2,454.0,115.63,17.01,3243.45,0,0,95350
6167,1,0,1,1,47,1,0,Fiber optic,1,0,0,1,Month-to-month,0,Electronic check,90.05,4137.2,0,57,20,38.25,3291,0,Modesto,1,1,Cable,37.621458000000004,-121.012295,1,90.05,1,3,None,47536,0,0,1,1,47,1,0.0,1797.75,0.0,4137.2,0,1,95351
6168,1,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.25,79.25,1,49,6,19.98,5533,1,Modesto,0,1,DSL,37.639029,-120.964772,0,82.42,0,0,Offer E,27135,0,1,0,1,1,5,0.0,19.98,0.0,79.25,0,1,95354
6169,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),44.9,44.9,1,30,65,41.78,2632,1,Modesto,0,0,DSL,37.672906,-120.94659399999999,0,46.696000000000005,0,0,Offer E,47613,0,1,0,0,1,5,0.0,41.78,0.0,44.9,0,0,95355
6170,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.4,19.4,0,49,0,2.85,5566,0,Modesto,0,0,NA,37.716186,-121.02583600000001,0,19.4,0,0,None,26055,0,0,0,0,1,2,0.0,2.85,0.0,19.4,0,0,95356
6171,0,1,1,1,59,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),88.75,5348.65,0,75,26,16.15,6492,0,Modesto,1,0,DSL,37.670526,-120.877572,1,88.75,1,3,None,13343,0,0,1,0,59,0,139.06,952.85,0.0,5348.65,0,1,95357
6172,1,0,1,0,10,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.1,659.65,1,42,21,22.03,2457,1,Modesto,0,1,Cable,37.612612,-121.10856799999999,1,72.904,0,1,None,30668,0,0,1,0,10,0,139.0,220.3,34.69,659.65,0,0,95358
6173,1,1,0,0,35,1,1,Fiber optic,1,0,0,1,Month-to-month,0,Credit card (automatic),91.0,3180.5,0,78,19,26.19,5527,0,Newman,0,1,DSL,37.343846,-121.039391,0,91.0,0,0,None,8504,0,1,0,0,35,3,604.0,916.65,0.0,3180.5,0,0,95360
6174,1,0,0,0,4,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,29.65,118.5,1,27,53,0.0,4207,1,Oakdale,1,1,Cable,37.785033,-120.776141,0,30.836,0,0,Offer E,25384,0,0,0,1,4,6,63.0,0.0,0.0,118.5,1,0,95361
6175,1,0,1,1,32,1,0,Fiber optic,1,1,0,1,One year,1,Electronic check,90.8,3023.85,0,29,69,36.65,2722,0,Patterson,0,1,Fiber Optic,37.410236,-121.32033700000001,1,90.8,3,6,None,15536,0,0,1,1,32,0,2086.0,1172.8,0.0,3023.85,1,0,95363
6176,1,0,0,0,43,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,77.85,3365.85,1,47,28,49.13,5107,1,Pinecrest,0,1,Cable,38.224869,-119.755729,0,80.964,0,0,Offer B,235,0,0,0,0,43,1,942.0,2112.59,0.0,3365.85,0,0,95364
6177,1,0,0,0,4,1,0,DSL,0,0,0,1,Month-to-month,0,Electronic check,54.3,195.3,1,64,21,40.15,5834,1,Planada,0,1,Fiber Optic,37.329725,-120.306399,0,56.472,0,0,Offer E,4150,0,0,0,1,4,2,0.0,160.6,0.0,195.3,0,1,95365
6178,0,1,1,0,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,18.95,1031.1,0,68,0,23.94,5548,0,Ripon,0,0,NA,37.750778000000004,-121.13238,1,18.95,0,3,None,12646,0,0,1,0,54,0,0.0,1292.76,0.0,1031.1,0,0,95366
6179,0,1,0,0,11,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),95.15,997.65,1,67,24,3.62,4074,1,Riverbank,0,0,Cable,37.734971,-120.95427099999999,0,98.956,0,0,None,16525,0,0,0,1,11,1,239.0,39.82,0.0,997.65,0,0,95367
6180,0,1,0,0,66,1,1,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),102.4,6471.85,0,68,20,10.45,4861,0,Salida,0,0,Cable,37.713152,-121.08738999999998,0,102.4,0,0,None,12466,0,0,0,1,66,1,0.0,689.6999999999998,0.0,6471.85,0,1,95368
6181,1,0,1,1,61,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,99.9,6241.35,0,62,58,34.54,5641,0,Snelling,1,1,Fiber Optic,37.521708000000004,-120.42684299999999,1,99.9,3,3,None,1158,0,1,1,1,61,1,3620.0,2106.94,0.0,6241.35,0,0,95369
6182,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),88.7,6501.35,0,64,19,28.63,4641,0,Sonora,1,1,DSL,37.982715999999996,-120.343732,1,88.7,2,1,Offer A,25340,1,1,1,1,72,1,1235.0,2061.36,0.0,6501.35,0,0,95370
6183,1,0,1,1,44,0,No phone service,DSL,0,0,1,1,One year,1,Electronic check,54.3,2317.1,0,25,69,0.0,3423,0,Soulsbyville,1,1,DSL,37.990574,-120.261821,1,54.3,1,1,None,1519,1,0,1,1,44,0,159.88,0.0,0.0,2317.1,1,1,95372
6184,1,0,0,0,41,1,1,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),55.7,2237.55,0,40,3,6.6,5590,0,Stevinson,1,1,Fiber Optic,37.316807,-120.855753,0,55.7,0,0,None,1960,0,0,0,0,41,2,0.0,270.6,0.0,2237.55,0,1,95374
6185,1,0,1,0,50,1,1,Fiber optic,1,0,1,1,One year,1,Electronic check,103.95,5231.3,0,27,51,23.28,4363,0,Tracy,1,1,Fiber Optic,37.680968,-121.446049,1,103.95,0,0,None,69801,0,0,0,1,50,0,0.0,1164.0,0.0,5231.3,1,1,95376
6186,1,0,1,0,47,1,1,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),110.85,5275.8,1,42,19,19.02,3344,1,Tuolumne,1,1,DSL,37.939768,-120.188002,1,115.284,0,1,Offer B,3979,1,0,1,1,47,1,1002.0,893.9399999999998,4.93,5275.8,0,0,95379
6187,1,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.15,165.5,0,30,0,2.87,3899,0,Turlock,0,1,NA,37.474396,-120.87591699999999,1,20.15,3,1,Offer E,40545,0,0,1,0,8,1,0.0,22.96,0.0,165.5,0,0,95380
6188,1,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,358.5,0,61,0,22.97,4204,0,Turlock,0,1,NA,37.529656,-120.85435700000001,0,20.05,0,0,None,24708,0,0,0,0,18,2,0.0,413.46,0.0,358.5,0,0,95382
6189,1,0,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),91.95,6614.9,0,21,59,27.1,4403,0,Twain Harte,1,1,Fiber Optic,38.107440999999994,-120.230625,1,91.95,1,1,Offer A,4848,1,0,1,1,72,0,0.0,1951.2,0.0,6614.9,1,1,95383
6190,1,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,0,Electronic check,80.5,80.5,1,24,76,35.77,2734,1,Vernalis,0,1,Cable,37.609095,-121.26338100000001,0,83.72,0,0,None,274,0,2,0,1,1,4,0.0,35.77,0.0,80.5,1,0,95385
6191,0,1,0,0,42,1,1,DSL,0,0,0,0,Month-to-month,0,Electronic check,55.65,2421.75,0,66,30,27.0,5831,0,Waterford,1,0,Cable,37.669515999999994,-120.62696399999999,0,55.65,0,0,None,8308,0,0,0,0,42,0,0.0,1134.0,0.0,2421.75,0,1,95386
6192,0,1,0,0,18,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,74.7,1294.6,0,78,18,21.09,3896,0,Escondido,0,0,Fiber Optic,33.141265000000004,-116.967221,0,74.7,0,0,Offer D,48690,0,0,0,0,18,0,233.0,379.62,0.0,1294.6,0,0,92027
6193,0,0,0,1,13,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),104.15,1299.1,0,29,27,11.99,2810,0,Winton,1,0,Cable,37.421299,-120.59958700000001,0,104.15,2,0,Offer D,11463,0,0,0,1,13,0,35.08,155.87,2.76,1299.1,1,1,95388
6194,0,0,1,1,68,1,1,Fiber optic,0,1,0,0,One year,1,Bank transfer (automatic),83.65,5733.4,0,50,29,15.94,5958,0,Escondido,0,0,Fiber Optic,33.141265000000004,-116.967221,1,83.65,2,1,Offer A,48690,1,0,1,0,68,0,1663.0,1083.92,46.99,5733.4,0,0,92027
6195,1,0,0,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),72.2,305.55,1,20,78,29.98,5668,1,Santa Rosa,0,1,Cable,38.460516999999996,-122.79033500000001,0,75.08800000000002,0,0,Offer E,36125,0,1,0,1,4,5,23.83,119.92,0.0,305.55,1,1,95401
6196,1,0,0,0,69,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),110.05,7430.75,0,27,73,5.71,5798,0,Santa Rosa,1,1,DSL,38.488431,-122.752839,0,110.05,0,0,Offer A,40270,0,0,0,1,69,0,5424.0,393.99,23.16,7430.75,1,0,95403
6197,1,0,0,0,17,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,51.5,900.5,1,36,2,46.6,5659,1,Santa Rosa,0,1,DSL,38.526941,-122.709096,0,53.56,0,0,Offer D,35057,1,1,0,0,17,4,0.0,792.2,35.34,900.5,0,1,95404
6198,1,0,1,1,25,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.5,630.6,0,31,0,23.69,5230,0,Santa Rosa,0,1,NA,38.439696000000005,-122.66881699999999,1,25.5,3,1,None,22250,0,0,1,0,25,2,0.0,592.25,44.42,630.6,0,0,95405
6199,1,1,0,0,43,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,89.55,3856.75,1,74,7,39.12,3802,1,Santa Rosa,0,1,Cable,38.394090999999996,-122.739814,0,93.132,0,0,None,30876,0,1,0,1,43,1,270.0,1682.16,0.0,3856.75,0,0,95407
6200,0,0,1,1,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.5,1222.65,0,19,0,9.51,4579,0,Santa Rosa,0,0,NA,38.468893,-122.58053899999999,1,19.5,2,1,None,25718,0,0,1,0,59,0,0.0,561.09,0.0,1222.65,1,0,95409
6201,0,1,0,0,5,1,0,Fiber optic,1,1,0,0,Month-to-month,0,Electronic check,80.7,374.8,0,72,17,36.27,3468,0,Albion,0,0,DSL,39.225694,-123.717354,0,80.7,0,0,Offer E,1054,0,0,0,0,5,1,64.0,181.35,0.0,374.8,0,0,95410
6202,1,0,1,1,21,1,1,DSL,1,1,1,0,One year,0,Mailed check,77.5,1625,1,34,15,17.57,5353,1,Annapolis,0,1,Cable,38.731055,-123.316553,1,80.60000000000002,0,1,Offer D,747,1,0,1,0,21,1,244.0,368.97,18.39,1625.0,0,0,95412
6203,0,0,1,1,69,1,1,Fiber optic,1,1,1,0,One year,1,Credit card (automatic),105.1,7234.8,0,19,48,23.02,4686,0,Boonville,1,0,Fiber Optic,39.025867,-123.38154399999999,1,105.1,3,1,Offer A,1374,1,0,1,0,69,0,3473.0,1588.38,0.0,7234.8,1,0,95415
6204,1,0,0,0,13,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),25.15,331.85,0,37,16,0.0,4943,0,Branscomb,0,1,DSL,39.710591,-123.682799,0,25.15,0,0,Offer D,176,0,0,0,0,13,2,0.0,0.0,48.59,331.85,0,1,95417
6205,1,0,1,0,42,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),95.25,3959.35,1,37,32,18.26,2075,1,Caspar,1,1,Cable,39.361283,-123.784599,1,99.06,0,1,Offer B,333,0,0,1,0,42,4,1267.0,766.9200000000002,27.3,3959.35,0,0,95420
6206,1,0,1,0,52,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),95.65,5088.4,0,27,85,8.94,4465,0,Cazadero,0,1,DSL,38.578807,-123.19338,1,95.65,0,1,None,1575,1,0,1,1,52,0,432.51,464.88,11.8,5088.4,1,1,95421
6207,1,1,0,0,46,1,0,Fiber optic,1,0,0,1,Month-to-month,0,Electronic check,85.0,3969.4,1,77,32,36.78,2097,1,Clearlake,0,1,Fiber Optic,38.965804,-122.63177900000001,0,88.4,0,0,None,13485,0,0,0,1,46,5,1270.0,1691.88,0.0,3969.4,0,0,95422
6208,1,0,1,0,61,1,1,DSL,1,1,0,1,Two year,1,Bank transfer (automatic),80.8,4860.85,0,53,20,43.48,4302,0,Clearlake Oaks,1,1,DSL,39.07116,-122.598542,1,80.8,0,1,None,3684,1,0,1,1,61,3,972.0,2652.28,17.17,4860.85,0,0,95423
6209,1,0,0,0,29,0,No phone service,DSL,0,0,0,0,One year,1,Mailed check,24.85,788.05,0,19,59,0.0,4161,0,Cloverdale,0,1,Fiber Optic,38.801936,-122.93893500000001,0,24.85,0,0,None,9210,0,0,0,0,29,1,46.49,0.0,0.0,788.05,1,1,95425
6210,0,0,0,1,25,1,0,DSL,0,1,0,0,One year,1,Credit card (automatic),54.75,1266.35,0,37,27,39.9,5136,0,Cobb,0,0,Cable,38.838088,-122.73203000000001,0,54.75,1,0,Offer C,1591,1,1,0,0,25,3,34.19,997.5,15.76,1266.35,0,1,95426
6211,0,0,1,1,5,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.75,470.95,1,38,24,1.12,3608,1,Comptche,0,0,Cable,39.239818,-123.565432,1,89.18,0,1,Offer E,371,1,0,1,0,5,5,113.0,5.6000000000000005,44.16,470.95,0,0,95427
6212,1,0,0,0,15,0,No phone service,DSL,0,0,1,1,One year,0,Electronic check,50.75,688.2,0,52,14,0.0,5091,0,Covelo,1,1,Fiber Optic,39.83307,-123.17876499999998,0,50.75,0,0,Offer D,2296,0,0,0,1,15,1,0.0,0.0,32.55,688.2,0,1,95428
6213,0,0,1,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.15,387.7,0,48,0,31.85,4246,0,Dos Rios,0,0,NA,39.756049,-123.358701,1,20.15,3,1,Offer D,91,0,0,1,0,19,0,0.0,605.15,2.97,387.7,0,0,95429
6214,1,0,0,0,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.05,845.25,0,28,0,47.53,2798,0,Duncans Mills,0,1,NA,38.445603000000006,-123.06375600000001,0,20.05,0,0,None,187,0,0,0,0,44,0,0.0,2091.32,15.31,845.25,1,0,95430
6215,0,1,0,0,6,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,98.25,560.6,1,79,32,47.35,3330,1,Lakewood,0,0,Cable,33.840524,-118.148403,0,102.18,0,0,None,30173,0,0,0,1,6,3,179.0,284.1,0.0,560.6,0,0,90712
6216,1,0,1,1,58,1,1,DSL,1,1,0,0,Two year,0,Credit card (automatic),71.6,4230.25,0,44,25,40.57,4747,0,Elk,1,1,Cable,39.108252,-123.645121,1,71.6,3,1,None,383,1,0,1,0,58,3,1058.0,2353.06,45.54,4230.25,0,0,95432
6217,1,0,1,1,62,1,0,Fiber optic,1,1,0,0,One year,1,Credit card (automatic),81.45,4983.05,0,27,41,39.67,5179,0,Forestville,0,1,Fiber Optic,38.499302,-122.92443999999999,1,81.45,3,1,None,6216,0,0,1,0,62,1,2043.0,2459.54,14.15,4983.05,1,0,95436
6218,0,0,1,1,70,0,No phone service,DSL,0,1,1,1,One year,1,Bank transfer (automatic),58.4,4113.15,0,52,19,0.0,4117,0,Fort Bragg,1,0,DSL,39.455555,-123.68397900000001,1,58.4,2,1,Offer A,14417,1,0,1,1,70,2,781.0,0.0,32.53,4113.15,0,0,95437
6219,0,1,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,25.7,25.7,1,68,10,0.0,4095,1,Fulton,0,0,Fiber Optic,38.493888,-122.77714099999999,0,26.728,0,0,None,476,0,0,0,0,1,3,0.0,0.0,0.0,25.7,0,0,95439
6220,1,0,1,1,10,0,No phone service,DSL,1,1,0,1,Two year,0,Credit card (automatic),53.7,521,0,49,24,0.0,5671,0,Geyserville,1,1,Fiber Optic,38.731771,-123.064272,1,53.7,2,2,Offer D,2349,1,0,1,1,10,1,0.0,0.0,22.97,521.0,0,1,95441
6221,1,0,0,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),19.6,471.85,0,64,0,37.7,3722,0,Glen Ellen,0,1,NA,38.368744,-122.52264199999999,0,19.6,0,0,Offer C,4101,0,0,0,0,26,3,0.0,980.2,21.25,471.85,0,0,95442
6222,1,0,0,0,66,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Credit card (automatic),89.4,5976.9,0,55,8,48.78,4889,0,Glenhaven,0,1,Fiber Optic,39.045246,-122.743181,0,89.4,0,0,Offer A,175,0,1,0,1,66,1,47.82,3219.48,36.02,5976.9,0,1,95443
6223,0,0,1,1,7,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.0,506.9,1,25,80,8.95,5672,1,Graton,0,0,Fiber Optic,38.434362,-122.86891000000001,1,71.76,0,1,Offer E,390,0,2,1,1,7,2,406.0,62.64999999999999,0.0,506.9,1,0,95444
6224,1,0,1,1,51,1,1,Fiber optic,0,1,0,0,One year,0,Bank transfer (automatic),84.2,4299.75,0,36,51,9.5,4952,0,Gualala,0,1,Fiber Optic,38.848082,-123.50608000000001,1,84.2,3,6,None,1916,1,0,1,0,51,1,0.0,484.5,39.68,4299.75,0,1,95445
6225,1,0,1,1,72,1,1,Fiber optic,1,1,1,0,Two year,1,Credit card (automatic),106.1,7548.6,0,31,24,7.16,4890,0,Guerneville,1,1,Cable,38.52576,-123.013347,1,106.1,1,9,Offer A,4913,1,0,1,0,72,3,181.17,515.52,23.39,7548.6,0,1,95446
6226,1,0,0,0,65,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.75,1654.75,0,56,0,4.9,5707,0,Healdsburg,0,1,NA,38.618347,-122.908422,0,25.75,0,0,None,17979,0,0,0,0,65,1,0.0,318.5,41.74,1654.75,0,0,95448
6227,1,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),46.05,80.35,1,27,57,29.69,4662,1,Hopland,0,1,DSL,38.937059999999995,-123.11811100000001,0,47.892,0,0,Offer E,1373,0,0,0,1,2,2,46.0,59.38,0.0,80.35,1,0,95449
6228,1,0,0,1,70,1,1,DSL,1,1,0,0,One year,0,Bank transfer (automatic),64.95,4551.5,0,31,19,26.62,5392,0,Jenner,0,1,Fiber Optic,38.505995,-123.18701899999999,0,64.95,1,0,None,438,1,1,0,0,70,1,865.0,1863.4,20.87,4551.5,0,0,95450
6229,1,0,1,0,72,1,1,DSL,0,1,1,1,Two year,1,Credit card (automatic),85.45,6227.5,0,39,16,31.15,5641,0,Kelseyville,1,1,Fiber Optic,38.93496,-122.792243,1,85.45,0,10,None,9902,1,1,1,1,72,1,0.0,2242.8,0.0,6227.5,0,1,95451
6230,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,20.05,0,61,0,16.02,5811,0,Kenwood,0,0,NA,38.419525,-122.52158500000002,1,20.05,3,3,None,1653,0,0,1,0,1,0,0.0,16.02,0.0,20.05,0,0,95452
6231,0,1,1,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Mailed check,76.4,76.4,1,76,7,41.16,2426,1,Lakeport,0,0,DSL,39.080469,-122.955176,1,79.456,0,6,None,11180,0,0,1,0,1,5,0.0,41.16,0.0,76.4,0,0,95453
6232,0,0,0,0,5,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.5,514,1,54,32,28.2,5180,1,Laytonville,1,0,Cable,39.806141,-123.531098,0,104.52,0,0,None,2706,0,1,0,1,5,2,0.0,141.0,0.0,514.0,0,1,95454
6233,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.7,57.5,0,27,0,38.41,2011,0,Little River,0,1,NA,39.245911,-123.77214,0,20.7,0,0,Offer E,882,0,0,0,0,3,0,0.0,115.23,0.0,57.5,1,0,95456
6234,1,0,0,0,58,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.3,1474.35,0,39,0,48.78,4477,0,Lower Lake,0,1,NA,38.925545,-122.54908300000001,0,25.3,0,0,None,2644,0,0,0,0,58,2,0.0,2829.24,0.0,1474.35,0,0,95457
6235,1,1,1,1,22,0,No phone service,DSL,1,0,0,1,Month-to-month,0,Mailed check,40.05,880.2,1,80,20,0.0,2061,1,Lucerne,0,1,Cable,39.141934,-122.770679,1,41.652,2,5,None,3002,0,0,1,0,22,0,176.0,0.0,0.0,880.2,0,0,95458
6236,1,1,1,0,33,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),100.6,3270.25,0,79,22,44.1,3669,0,Manchester,0,1,Fiber Optic,38.966713,-123.58641200000001,1,100.6,0,6,None,586,0,0,1,0,33,1,71.95,1455.3,0.0,3270.25,0,1,95459
6237,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.95,69.95,1,48,18,27.58,5066,1,Mendocino,0,1,Cable,39.305545,-123.743697,0,72.748,0,0,Offer E,2229,0,0,0,0,1,4,0.0,27.58,0.0,69.95,0,0,95460
6238,1,1,1,0,54,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),74.0,3919.15,0,73,5,35.16,4991,0,Middletown,0,1,DSL,38.787446,-122.58675,1,74.0,0,10,None,7789,0,0,1,0,54,2,0.0,1898.64,0.0,3919.15,0,1,95461
6239,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,99.4,7285.7,0,21,48,34.95,6022,0,Monte Rio,0,1,Fiber Optic,38.471049,-123.015549,1,99.4,0,7,None,1537,0,0,1,1,72,3,3497.0,2516.4,0.0,7285.7,1,0,95462
6240,1,0,0,1,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.3,93.3,1,59,33,7.99,2578,1,Navarro,0,1,DSL,39.182916,-123.552571,0,97.03200000000001,0,0,Offer E,148,0,0,0,1,1,2,0.0,7.99,0.0,93.3,0,0,95463
6241,1,0,0,0,3,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,49.15,169.05,1,47,32,40.79,5598,1,Nice,1,1,Cable,39.12334,-122.83819799999999,0,51.11600000000001,0,0,Offer E,2223,0,1,0,0,3,6,54.0,122.37,0.0,169.05,0,0,95464
6242,0,0,1,1,72,1,1,Fiber optic,1,1,0,1,Two year,0,Credit card (automatic),107.45,7658.3,0,35,19,17.89,4505,0,Occidental,1,0,DSL,38.415003000000006,-122.998726,1,107.45,2,1,None,1880,1,1,1,1,72,1,1455.0,1288.08,0.0,7658.3,0,0,95465
6243,0,0,1,1,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),83.6,5959.3,0,36,22,12.84,4116,0,Philo,1,0,DSL,39.094102,-123.500853,1,83.6,1,4,None,1113,0,1,1,1,72,2,0.0,924.48,0.0,5959.3,0,1,95466
6244,1,1,1,0,54,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Credit card (automatic),99.05,5295.7,0,67,13,38.48,4011,0,Point Arena,1,1,Cable,38.911299,-123.60958799999999,1,99.05,0,0,None,1352,0,0,0,0,54,0,0.0,2077.92,0.0,5295.7,0,1,95468
6245,0,0,1,0,59,1,1,DSL,0,1,1,1,One year,1,Electronic check,80.1,4693.2,0,34,13,20.27,4093,0,Potter Valley,0,0,Fiber Optic,39.408634,-123.04551599999999,1,80.1,0,7,None,1884,1,0,1,1,59,0,61.01,1195.93,0.0,4693.2,0,1,95469
6246,1,0,0,0,54,1,0,DSL,1,1,1,0,Two year,1,Bank transfer (automatic),65.3,3512.9,0,47,16,18.74,4556,0,Redwood Valley,0,1,Fiber Optic,39.298065,-123.25211000000002,0,65.3,0,0,None,5995,0,1,0,0,54,2,0.0,1011.96,0.0,3512.9,0,1,95470
6247,1,0,0,0,60,1,1,Fiber optic,0,0,1,0,Two year,1,Electronic check,89.55,5231.2,0,34,10,7.1,5874,0,Rio Nido,1,1,Fiber Optic,38.522328,-122.97932,0,89.55,0,0,None,298,0,0,0,0,60,2,523.0,426.0,0.0,5231.2,0,0,95471
6248,0,0,1,0,60,0,No phone service,DSL,0,1,1,1,Two year,0,Credit card (automatic),60.8,3603.45,0,19,69,0.0,5784,0,Sebastopol,1,0,Cable,38.398815,-122.861923,1,60.8,0,5,None,31266,1,0,1,1,60,0,0.0,0.0,0.0,3603.45,1,1,95472
6249,1,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,74.5,217.45,0,39,14,6.97,5203,0,Sonoma,0,1,Cable,38.25485,-122.461799,0,74.5,0,0,None,34314,0,0,0,0,3,1,0.0,20.91,0.0,217.45,0,1,95476
6250,0,0,1,0,69,1,1,Fiber optic,1,0,1,1,Two year,0,Bank transfer (automatic),99.15,6875.35,0,52,19,45.35,5031,0,Ukiah,0,0,Cable,39.134075,-123.23422,1,99.15,0,6,None,30988,0,0,1,1,69,2,1306.0,3129.15,0.0,6875.35,0,0,95482
6251,0,0,1,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Electronic check,19.25,19.25,0,29,0,25.1,2053,0,Upper Lake,0,0,NA,39.220368,-122.907693,1,19.25,5,9,Offer E,2344,0,0,1,0,1,0,0.0,25.1,0.0,19.25,1,0,95485
6252,1,0,1,1,50,0,No phone service,DSL,1,0,1,0,Month-to-month,1,Credit card (automatic),39.45,2021.35,0,44,23,0.0,6018,0,Westport,0,1,Fiber Optic,39.724433000000005,-123.767578,1,39.45,3,10,None,309,0,0,1,0,50,0,0.0,0.0,0.0,2021.35,0,1,95488
6253,0,0,0,0,56,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),44.85,2564.95,0,58,23,0.0,4021,0,Willits,0,0,Fiber Optic,39.492046,-123.375818,0,44.85,0,0,None,13472,0,0,0,1,56,0,58.99,0.0,0.0,2564.95,0,1,95490
6254,0,0,1,0,60,1,0,Fiber optic,1,0,1,1,Two year,1,Electronic check,97.2,5611.75,0,59,13,32.5,4905,0,Windsor,0,0,Fiber Optic,38.527297,-122.81004399999999,1,97.2,0,6,None,23701,1,0,1,1,60,1,0.0,1950.0,0.0,5611.75,0,1,95492
6255,1,1,1,0,69,1,1,Fiber optic,1,0,1,1,One year,1,Mailed check,110.55,7610.1,0,73,14,8.3,4887,0,Witter Springs,1,1,DSL,39.222322999999996,-122.98548799999999,1,110.55,0,2,None,240,1,0,1,0,69,1,0.0,572.7,0.0,7610.1,0,1,95493
6256,0,0,0,0,1,0,No phone service,DSL,0,0,0,1,Month-to-month,0,Mailed check,35.05,35.05,1,62,24,0.0,3706,1,Yorkville,0,0,Cable,38.888351,-123.23964699999999,0,36.452,0,0,Offer E,335,0,2,0,1,1,2,0.0,0.0,0.0,35.05,0,0,95494
6257,0,1,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,73.0,73,1,72,6,20.55,4116,1,The Sea Ranch,0,0,Cable,38.696659000000004,-123.43686100000001,0,75.92,0,0,None,752,0,1,0,0,1,3,0.0,20.55,0.0,73.0,0,0,95497
6258,0,0,1,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.9,45.75,0,55,0,41.36,3716,0,Eureka,0,0,NA,40.796621,-124.15428,1,19.9,0,4,Offer E,23224,0,0,1,0,3,2,0.0,124.08,0.0,45.75,0,0,95501
6259,1,0,1,1,60,1,0,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),76.95,4543.95,0,39,21,27.2,5053,0,Eureka,0,1,DSL,40.737431,-124.108897,1,76.95,3,7,None,23570,1,0,1,1,60,0,954.0,1632.0,0.0,4543.95,0,0,95503
6260,0,0,0,0,13,0,No phone service,DSL,0,0,0,0,Two year,0,Mailed check,35.4,450.4,0,58,13,0.0,3239,0,Alderpoint,1,0,Fiber Optic,40.166028000000004,-123.584144,0,35.4,0,0,Offer D,261,1,0,0,0,13,0,59.0,0.0,0.0,450.4,0,0,95511
6261,1,0,1,1,62,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.45,1297.35,0,45,0,1.87,5746,0,Blocksburg,0,1,NA,40.309088,-123.668201,1,20.45,2,2,None,199,0,0,1,0,62,0,0.0,115.94,0.0,1297.35,0,0,95514
6262,0,0,0,0,45,1,1,Fiber optic,1,1,0,1,One year,0,Bank transfer (automatic),96.75,4442.75,0,58,30,1.57,3682,0,Mckinleyville,0,0,Fiber Optic,40.965011,-124.01525500000001,0,96.75,0,0,None,15921,0,1,0,1,45,1,133.28,70.65,0.0,4442.75,0,1,95519
6263,0,0,0,0,25,0,No phone service,DSL,0,0,1,1,One year,0,Electronic check,54.2,1423.15,0,37,29,0.0,4458,0,Arcata,1,0,Cable,40.839958,-124.00375700000001,0,54.2,0,0,Offer C,19596,1,1,0,1,25,2,41.27,0.0,0.0,1423.15,0,1,95521
6264,1,0,0,0,44,1,0,Fiber optic,0,0,1,1,Two year,0,Bank transfer (automatic),100.1,4378.35,0,30,59,48.95,4025,0,Bayside,1,1,DSL,40.825486,-124.049485,0,100.1,0,0,Offer B,1689,1,0,0,1,44,2,2583.0,2153.8,0.0,4378.35,0,0,95524
6265,0,0,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.25,74.2,0,34,26,39.5,5441,0,Blue Lake,0,0,DSL,40.94338,-123.831799,0,45.25,0,0,Offer E,1584,0,0,0,0,2,2,0.0,79.0,0.0,74.2,0,1,95525
6266,1,1,0,0,33,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),83.85,2716.3,1,78,2,38.53,2583,1,Bridgeville,1,1,Fiber Optic,40.372532,-123.525626,0,87.204,0,0,None,695,0,0,0,0,33,4,54.0,1271.49,0.0,2716.3,0,0,95526
6267,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.1,70.1,1,43,28,17.37,3706,1,Burnt Ranch,0,0,Fiber Optic,40.854512,-123.450097,0,72.904,0,0,None,485,0,1,0,0,1,4,0.0,17.37,0.0,70.1,0,0,95527
6268,0,0,0,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.85,450.65,0,50,0,10.25,3171,0,Carlotta,0,0,NA,40.497283,-123.93037,0,20.85,0,0,Offer D,1072,0,0,0,0,22,0,0.0,225.5,0.0,450.65,0,0,95528
6269,0,0,0,0,35,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,33.45,1175.85,0,59,12,0.0,2553,0,Fallbrook,1,0,Cable,33.362575,-117.299644,0,33.45,0,0,Offer C,42239,1,0,0,0,35,1,14.11,0.0,0.0,1175.85,0,1,92028
6270,0,0,1,1,29,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.2,558.8,0,40,0,34.44,2784,0,Ferndale,0,0,NA,40.4785,-124.301372,1,20.2,1,5,Offer C,2965,0,0,1,0,29,0,0.0,998.76,0.0,558.8,0,0,95536
6271,1,1,1,0,27,1,1,Fiber optic,1,0,0,0,One year,1,Electronic check,85.9,2220.1,0,72,14,41.11,5755,0,Fields Landing,1,1,DSL,40.726949,-124.217378,1,85.9,0,7,None,228,0,0,1,0,27,0,0.0,1109.97,0.0,2220.1,0,1,95537
6272,1,0,0,1,54,1,0,DSL,0,1,0,0,One year,1,Electronic check,61.0,3283.05,0,20,59,4.16,5594,0,Fortuna,1,1,Fiber Optic,40.584990999999995,-124.121504,0,61.0,2,0,Offer B,12241,1,0,0,0,54,0,1937.0,224.64,0.0,3283.05,1,0,95540
6273,0,1,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.65,142.35,1,67,28,12.52,2189,1,Garberville,0,0,DSL,40.057784000000005,-123.679461,0,73.47600000000001,0,0,None,2423,0,1,0,0,2,5,40.0,25.04,0.0,142.35,0,0,95542
6274,1,0,0,0,57,1,1,Fiber optic,0,0,1,0,One year,1,Electronic check,86.9,4939.25,0,45,26,36.08,6109,0,Gasquet,0,1,DSL,41.867908,-123.79414399999999,0,86.9,0,0,Offer B,532,0,0,0,0,57,1,0.0,2056.56,0.0,4939.25,0,1,95543
6275,1,0,0,0,62,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),69.4,4237.5,0,55,12,41.13,6469,0,Honeydew,1,1,Fiber Optic,40.342928,-124.06332900000001,0,69.4,0,0,Offer B,82,1,2,0,0,62,1,508.0,2550.06,0.0,4237.5,0,0,95545
6276,0,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),20.35,335.95,0,44,0,46.64,3205,0,Hoopa,0,0,NA,41.163637,-123.70484099999999,1,20.35,3,10,Offer D,3041,0,0,1,0,15,2,0.0,699.6,0.0,335.95,0,0,95546
6277,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,33.2,1,62,0,32.03,5627,1,Hydesville,0,1,NA,40.557314,-124.08166200000001,0,20.35,0,0,None,1201,0,1,0,0,2,4,0.0,64.06,0.0,33.2,0,0,95547
6278,0,0,1,0,70,1,1,Fiber optic,0,0,1,1,Two year,1,Bank transfer (automatic),104.3,7188.5,0,50,30,5.46,5583,0,Klamath,1,0,DSL,41.572813000000004,-124.03501100000001,1,104.3,0,9,None,1215,1,0,1,1,70,0,0.0,382.2,0.0,7188.5,0,1,95548
6279,0,0,1,1,21,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.95,926.25,0,33,17,38.95,3752,0,Kneeland,0,0,Fiber Optic,40.664483000000004,-123.865325,1,44.95,2,6,Offer D,264,0,1,1,0,21,1,0.0,817.95,0.0,926.25,0,1,95549
6280,0,0,0,1,23,1,0,DSL,0,0,0,0,One year,1,Electronic check,49.45,1119.35,0,61,53,25.85,5237,0,Korbel,0,0,Fiber Optic,40.7666,-123.80458,0,49.45,3,0,Offer D,155,1,0,0,0,23,0,0.0,594.5500000000002,0.0,1119.35,0,1,95550
6281,1,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.6,116.6,0,24,0,12.17,4439,0,Loleta,0,1,NA,40.665952000000004,-124.240051,0,20.6,0,0,Offer E,1447,0,0,0,0,6,0,0.0,73.02,0.0,116.6,1,0,95551
6282,1,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.55,68.8,0,53,0,29.09,5573,0,Mad River,0,1,NA,40.390301,-123.412327,1,19.55,3,0,Offer E,265,0,0,0,0,4,1,0.0,116.36,0.0,68.8,0,0,95552
6283,0,0,0,0,3,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Credit card (automatic),99.0,287.4,1,29,65,33.39,5236,1,Miranda,1,0,Cable,40.210895,-123.86,0,102.96,0,0,None,867,0,1,0,1,3,2,187.0,100.17,0.0,287.4,1,0,95553
6284,0,0,0,0,23,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,93.5,2341.55,0,46,23,18.12,4861,0,Myers Flat,0,0,Fiber Optic,40.267158,-123.80591299999999,0,93.5,0,0,Offer D,644,0,0,0,1,23,1,53.86,416.7600000000001,0.0,2341.55,0,1,95554
6285,1,0,0,0,26,0,No phone service,DSL,1,0,1,1,One year,0,Credit card (automatic),54.55,1362.85,0,22,82,0.0,4296,0,Orick,0,1,Fiber Optic,41.336354,-124.044354,0,54.55,0,0,Offer C,494,1,0,0,1,26,1,0.0,0.0,0.0,1362.85,1,1,95555
6286,0,0,0,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,163.6,0,24,0,15.66,2675,0,Orleans,0,0,NA,41.269521000000005,-123.546958,0,20.05,2,0,Offer E,574,0,0,0,0,8,1,0.0,125.28,0.0,163.6,1,0,95556
6287,1,0,0,0,26,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,83.95,2254.2,1,36,22,14.3,5869,1,Petrolia,0,1,Cable,40.274302,-124.210902,0,87.30799999999999,0,0,None,300,0,0,0,1,26,2,0.0,371.8,0.0,2254.2,0,1,95558
6288,1,0,0,0,2,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.45,145.15,0,20,85,28.61,2657,0,Phillipsville,0,1,Fiber Optic,40.184094,-123.74548700000001,0,79.45,0,0,Offer E,163,0,1,0,0,2,1,123.0,57.22,0.0,145.15,1,0,95559
6289,1,0,0,0,67,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),116.2,7752.3,1,25,78,33.88,4495,1,Redway,1,1,DSL,40.142256,-123.85292700000001,0,120.848,0,0,Offer A,1851,1,0,0,1,67,4,6047.0,2269.96,0.0,7752.3,1,0,95560
6290,0,0,1,0,71,1,1,Fiber optic,0,0,1,1,Two year,1,Bank transfer (automatic),93.7,6585.35,1,55,19,40.52,4296,1,Rio Dell,0,0,DSL,40.485849,-124.163234,1,97.448,0,2,Offer A,3284,0,0,1,1,71,2,0.0,2876.92,0.0,6585.35,0,1,95562
6291,0,0,0,0,59,1,1,DSL,1,1,0,1,One year,0,Credit card (automatic),79.85,4786.1,0,26,73,1.94,6041,0,Salyer,1,0,DSL,40.89866,-123.539754,0,79.85,0,0,Offer B,660,1,0,0,1,59,1,0.0,114.46,0.0,4786.1,1,1,95563
6292,1,0,1,1,39,1,1,Fiber optic,0,0,1,1,One year,0,Electronic check,100.0,3835.55,0,62,75,17.29,5434,0,Samoa,1,1,Cable,40.809636,-124.189977,1,100.0,3,9,Offer C,395,0,0,1,1,39,1,0.0,674.31,0.0,3835.55,0,1,95564
6293,1,0,0,1,21,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.6,397,0,45,0,27.6,2447,0,Scotia,0,1,NA,40.440636,-124.098739,0,19.6,2,0,Offer D,1125,0,0,0,0,21,0,0.0,579.6,0.0,397.0,0,0,95565
6294,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.7,19.7,1,42,0,1.91,5707,1,Smith River,0,1,NA,41.950683000000005,-124.097094,0,19.7,0,0,None,2020,0,0,0,0,1,2,0.0,1.91,0.0,19.7,0,0,95567
6295,0,0,1,1,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.2,1027.25,0,60,0,18.64,3828,0,Somes Bar,0,0,NA,41.444606,-123.47189499999999,1,20.2,2,6,Offer B,202,0,0,1,0,48,0,0.0,894.72,0.0,1027.25,0,0,95568
6296,0,1,1,0,31,0,No phone service,DSL,1,1,0,1,One year,1,Credit card (automatic),50.4,1580.1,0,72,21,0.0,2166,0,Redcrest,1,0,Cable,40.363446,-123.83504099999999,1,50.4,0,10,Offer C,400,0,0,1,0,31,0,332.0,0.0,0.0,1580.1,0,0,95569
6297,0,0,1,1,64,1,1,Fiber optic,1,1,1,1,One year,0,Electronic check,113.35,7222.75,0,63,19,6.83,4952,0,Trinidad,1,0,Fiber Optic,41.162295,-124.027381,1,113.35,1,1,Offer B,2369,1,0,1,1,64,0,0.0,437.12,0.0,7222.75,0,1,95570
6298,1,0,1,1,46,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.0,3769.7,0,43,16,5.52,3315,0,Weott,0,1,Cable,40.310119,-123.909449,1,80.0,1,1,Offer B,270,0,0,1,0,46,0,603.0,253.92,0.0,3769.7,0,0,95571
6299,0,0,0,0,52,1,1,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),80.95,4233.95,0,32,21,38.71,4924,0,Willow Creek,1,0,Fiber Optic,40.949011999999996,-123.655847,0,80.95,0,0,Offer B,1666,1,0,0,1,52,0,0.0,2012.92,0.0,4233.95,0,1,95573
6300,0,0,1,1,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,24.9,1680.25,0,54,0,17.43,5847,0,Leggett,0,0,NA,39.873371,-123.741474,1,24.9,1,4,None,321,0,0,1,0,67,0,0.0,1167.81,0.0,1680.25,0,0,95585
6301,0,1,0,0,67,1,1,DSL,0,1,0,0,Month-to-month,0,Electronic check,54.9,3725.5,0,68,28,48.43,4826,0,Piercy,0,0,Cable,39.955587,-123.681175,0,54.9,0,0,None,200,0,2,0,0,67,1,0.0,3244.81,0.0,3725.5,0,1,95587
6302,0,0,0,0,5,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.55,413.65,1,20,64,35.22,4600,1,Fallbrook,0,0,Cable,33.362575,-117.299644,0,78.572,0,0,None,42239,0,1,0,1,5,5,26.47,176.1,0.0,413.65,1,1,92028
6303,0,0,1,0,71,1,1,Fiber optic,0,1,1,1,Two year,0,Electronic check,109.25,7707.7,0,32,22,29.78,5044,0,Zenia,1,0,Fiber Optic,40.170357,-123.417298,1,109.25,0,7,None,259,1,0,1,1,71,0,169.57,2114.38,0.0,7707.7,0,1,95595
6304,0,0,0,0,9,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),77.65,714.15,1,40,25,22.88,3847,1,Amador City,0,0,DSL,38.431407,-120.8421,0,80.75600000000001,0,0,None,222,0,0,0,0,9,0,179.0,205.92,0.0,714.15,0,0,95601
6305,0,1,0,0,26,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Electronic check,95.0,2497.2,1,74,29,47.63,4232,1,Auburn,0,0,Cable,38.99003,-121.11440800000001,0,98.8,0,0,None,18197,0,0,0,0,26,6,0.0,1238.38,0.0,2497.2,0,1,95602
6306,1,0,0,0,71,1,1,Fiber optic,1,1,1,1,One year,1,Bank transfer (automatic),116.3,8309.55,0,22,48,2.88,4644,0,Auburn,1,1,DSL,38.912881,-121.08276599999999,0,116.3,0,0,None,24944,1,0,0,1,71,0,0.0,204.48,0.0,8309.55,1,1,95603
6307,0,0,0,0,32,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.9,601.55,0,35,0,15.53,4374,0,West Sacramento,0,0,NA,38.592745,-121.54003600000001,0,19.9,0,0,Offer C,12756,0,0,0,0,32,0,0.0,496.96,0.0,601.55,0,0,95605
6308,0,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.35,139.25,0,32,9,44.77,3430,0,Brooks,0,0,Fiber Optic,38.809804,-122.24138300000001,0,70.35,0,0,None,382,0,0,0,0,2,2,13.0,89.54,0.0,139.25,0,0,95606
6309,0,0,1,0,71,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.6,1888.25,0,48,0,11.18,5063,0,Capay,0,0,NA,38.681651,-122.130569,1,25.6,0,3,None,262,0,0,1,0,71,1,0.0,793.78,0.0,1888.25,0,0,95607
6310,0,0,0,0,60,0,No phone service,DSL,1,0,0,1,One year,1,Electronic check,44.45,2773.9,0,29,73,0.0,4928,0,Carmichael,1,0,DSL,38.626128,-121.328011,0,44.45,0,0,Offer B,58830,0,0,0,1,60,1,2025.0,0.0,0.0,2773.9,1,0,95608
6311,0,1,0,0,55,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,100.15,5409.75,0,75,3,29.6,5182,0,Citrus Heights,1,0,Fiber Optic,38.69508,-121.271616,0,100.15,0,0,None,43718,0,0,0,0,55,3,162.0,1628.0,0.0,5409.75,0,0,95610
6312,1,0,0,0,54,1,0,Fiber optic,1,1,1,1,One year,1,Credit card (automatic),105.4,5643.4,1,31,29,49.98,4406,1,Clarksburg,0,1,Cable,38.384648,-121.578701,0,109.616,0,0,Offer B,1417,1,4,0,1,54,2,1637.0,2698.92,0.0,5643.4,0,0,95612
6313,1,0,0,0,2,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.85,197.7,1,63,20,37.43,3790,1,Cool,1,1,Cable,38.880621999999995,-120.97386499999999,0,99.684,0,0,None,3674,0,1,0,1,2,4,40.0,74.86,0.0,197.7,0,0,95614
6314,0,0,0,0,6,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,73.85,401.3,0,45,9,27.69,4220,0,Courtland,0,0,Cable,38.311609000000004,-121.554034,0,73.85,0,0,None,699,0,0,0,0,6,2,0.0,166.14,0.0,401.3,0,1,95615
6315,0,0,1,1,48,1,0,DSL,1,1,0,1,Two year,1,Credit card (automatic),70.1,3238.4,0,56,57,4.45,5476,0,Davis,1,0,Fiber Optic,38.508734999999994,-121.67881299999999,1,70.1,3,1,Offer B,67411,0,0,1,1,48,2,1846.0,213.6,0.0,3238.4,0,0,95616
6316,1,0,1,1,63,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.25,1573.05,0,19,0,24.5,6245,0,Davis,0,1,NA,38.544002,-121.68555900000001,1,25.25,3,8,Offer B,648,0,0,1,0,63,0,0.0,1543.5,0.0,1573.05,1,0,95618
6317,1,0,0,0,1,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,79.15,79.15,1,64,26,24.48,4243,1,Diamond Springs,0,1,DSL,38.683605,-120.811852,0,82.316,0,0,None,4426,0,2,0,0,1,1,0.0,24.48,0.0,79.15,0,0,95619
6318,1,0,0,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),21.05,235.8,0,19,0,19.38,4001,0,Dixon,0,1,NA,38.392821000000005,-121.799917,0,21.05,2,0,Offer D,18529,0,0,0,0,12,1,0.0,232.56,0.0,235.8,1,0,95620
6319,1,1,1,0,54,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),24.95,1364.75,0,76,4,0.0,4691,0,Citrus Heights,0,1,Fiber Optic,38.69549,-121.307864,1,24.95,0,4,Offer B,41636,0,0,1,0,54,0,55.0,0.0,0.0,1364.75,0,0,95621
6320,0,0,1,1,30,1,0,DSL,0,0,1,0,One year,1,Electronic check,64.5,1985.15,0,56,18,36.74,2215,0,El Dorado,1,0,Fiber Optic,38.63153,-120.84260900000001,1,64.5,1,4,Offer C,4097,1,0,1,0,30,2,0.0,1102.2,0.0,1985.15,0,1,95623
6321,0,0,1,0,30,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.65,655.85,1,42,0,15.36,2486,1,Elk Grove,0,0,NA,38.434138,-121.30587,1,19.65,0,1,None,38534,0,1,1,0,30,2,0.0,460.8,0.0,655.85,0,0,95624
6322,0,0,0,0,4,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.0,303.15,1,61,30,27.57,2085,1,Elmira,0,0,Fiber Optic,38.349195,-121.902943,0,82.16,0,0,None,171,0,0,0,0,4,0,0.0,110.28,0.0,303.15,0,1,95625
6323,0,0,0,0,40,1,1,Fiber optic,0,0,1,1,One year,1,Credit card (automatic),105.95,4335.2,0,41,14,16.73,3784,0,Elverta,1,0,DSL,38.734997,-121.463719,0,105.95,0,0,Offer B,6197,1,0,0,1,40,2,0.0,669.2,0.0,4335.2,0,1,95626
6324,0,0,1,1,9,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.85,647.5,0,39,20,8.1,4843,0,Esparto,0,0,Fiber Optic,38.834469,-122.12719299999999,1,75.85,1,10,None,2756,1,0,1,0,9,1,0.0,72.89999999999998,0.0,647.5,0,1,95627
6325,0,0,1,1,17,1,0,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,91.85,1574.45,1,30,56,41.95,5643,1,Fair Oaks,0,0,DSL,38.652065,-121.25441000000001,1,95.524,0,1,Offer D,40750,1,0,1,0,17,2,882.0,713.1500000000002,0.0,1574.45,0,0,95628
6326,0,0,0,0,62,0,No phone service,DSL,0,1,0,1,Two year,1,Credit card (automatic),43.6,2748.7,0,38,30,0.0,4507,0,Fiddletown,1,0,Fiber Optic,38.513484000000005,-120.704613,0,43.6,0,0,Offer B,850,0,0,0,1,62,4,0.0,0.0,0.0,2748.7,0,1,95629
6327,1,0,0,0,28,1,0,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),91.25,2483.65,0,50,12,13.69,2886,0,Folsom,0,1,Cable,38.672638,-121.147403,0,91.25,0,0,Offer C,51855,1,0,0,0,28,0,0.0,383.32,0.0,2483.65,0,1,95630
6328,0,0,0,0,70,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),89.75,6367.2,0,64,7,29.53,5150,0,Foresthill,1,0,Fiber Optic,39.031876000000004,-120.81114099999999,0,89.75,0,0,None,5714,1,0,0,1,70,2,0.0,2067.1,0.0,6367.2,0,1,95631
6329,0,0,0,0,46,1,0,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),104.4,4904.2,0,20,82,5.86,4190,0,Galt,1,0,Fiber Optic,38.274451,-121.259201,0,104.4,0,0,Offer B,24194,1,1,0,1,46,2,0.0,269.56,0.0,4904.2,1,1,95632
6330,0,0,1,0,23,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Mailed check,90.15,2044.95,0,33,15,22.17,5110,0,Garden Valley,1,0,DSL,38.852544,-120.83766899999999,1,90.15,0,2,Offer D,2536,0,0,1,1,23,0,30.67,509.91,0.0,2044.95,0,1,95633
6331,1,0,1,1,47,0,No phone service,DSL,1,0,0,0,One year,0,Electronic check,40.3,1794.8,0,27,47,0.0,5040,0,Georgetown,1,1,DSL,38.9386,-120.78551399999999,1,40.3,1,7,Offer B,2723,1,0,1,0,47,2,0.0,0.0,0.0,1794.8,1,1,95634
6332,1,0,1,1,68,1,0,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),105.25,7173.15,0,41,19,31.4,5795,0,Greenwood,1,1,Fiber Optic,38.921333000000004,-120.897718,1,105.25,2,3,None,1140,0,0,1,1,68,1,0.0,2135.2,0.0,7173.15,0,1,95635
6333,0,1,0,0,60,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,106.0,6441.4,1,68,19,34.39,5507,1,Grizzly Flats,1,0,Cable,38.636102,-120.522149,0,110.24,0,0,None,659,1,0,0,0,60,3,1224.0,2063.4,0.0,6441.4,0,0,95636
6334,0,0,0,1,67,1,1,Fiber optic,0,1,1,1,Two year,1,Electronic check,104.0,7039.05,0,28,59,12.54,4741,0,Guinda,0,0,Fiber Optic,38.830739,-122.196202,0,104.0,1,0,None,228,1,0,0,1,67,1,0.0,840.18,0.0,7039.05,1,1,95637
6335,0,0,0,0,14,1,0,DSL,0,0,1,1,Month-to-month,1,Electronic check,69.65,921.4,0,52,29,37.01,5351,0,Herald,0,0,DSL,38.313447,-121.12388600000001,0,69.65,0,0,Offer D,1745,1,2,0,1,14,3,267.0,518.14,0.0,921.4,0,0,95638
6336,1,0,1,1,57,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.3,4018.35,0,59,22,49.95,4133,0,Hood,0,1,DSL,38.375325,-121.507935,1,74.3,2,4,Offer B,213,0,0,1,0,57,1,884.0,2847.15,0.0,4018.35,0,0,95639
6337,0,0,1,1,55,1,1,Fiber optic,1,0,1,1,One year,0,Mailed check,100.9,5448.6,0,34,18,41.18,6153,0,Ione,0,0,Fiber Optic,38.33788,-120.954202,1,100.9,1,6,Offer B,9752,0,0,1,1,55,1,981.0,2264.9,0.0,5448.6,0,0,95640
6338,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.25,20.25,0,25,0,42.96,4769,0,Isleton,0,1,NA,38.154823,-121.601358,0,20.25,0,0,None,2010,0,0,0,0,1,2,0.0,42.96,0.0,20.25,1,0,95641
6339,1,0,0,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,49.9,49.9,1,34,19,39.6,3113,1,Jackson,0,1,DSL,38.336216,-120.76901000000001,0,51.896,1,0,None,6202,1,0,0,0,1,3,0.0,39.6,0.0,49.9,0,0,95642
6340,1,0,0,0,23,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),96.9,2085.45,0,61,6,8.5,3875,0,Knights Landing,1,1,Fiber Optic,38.875508,-121.76586599999999,0,96.9,0,0,Offer D,1793,1,0,0,0,23,0,0.0,195.5,0.0,2085.45,0,1,95645
6341,0,0,0,0,13,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,100.35,1358.85,1,54,29,6.78,2008,1,Kirkwood,0,0,Fiber Optic,38.631489,-120.01516699999999,0,104.36399999999999,0,0,Offer D,129,0,1,0,1,13,4,394.0,88.14,34.09,1358.85,0,0,95646
6342,1,0,1,0,47,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.1,5135.15,0,61,21,48.69,3142,0,Lincoln,1,1,DSL,38.922812,-121.312005,1,104.1,0,2,Offer B,15286,0,0,1,1,47,2,0.0,2288.43,0.0,5135.15,0,1,95648
6343,1,0,0,0,38,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,730.1,0,38,0,22.23,2907,0,Loomis,0,1,NA,38.809175,-121.171375,0,20.1,0,0,None,11191,0,1,0,0,38,3,0.0,844.74,0.0,730.1,0,0,95650
6344,0,1,1,0,38,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.95,2869.85,1,66,33,15.78,5165,1,Lotus,0,0,DSL,38.815515000000005,-120.916997,1,77.94800000000002,0,5,None,485,0,3,1,0,38,1,947.0,599.64,0.0,2869.85,0,0,95651
6345,0,1,0,0,2,1,1,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),56.55,118.25,0,68,25,31.74,2069,0,Madison,0,0,Fiber Optic,38.674276,-121.96186599999999,0,56.55,0,0,Offer E,844,0,0,0,0,2,0,0.0,63.48,0.0,118.25,0,1,95653
6346,1,1,1,1,1,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),49.25,49.25,1,71,21,8.38,4478,1,Mather,0,1,Fiber Optic,38.549822,-121.266725,1,51.22,1,3,None,929,1,1,1,0,1,4,0.0,8.38,0.0,49.25,0,0,95655
6347,1,0,1,0,15,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),68.6,1108.6,0,54,10,24.17,3351,0,Newcastle,0,1,Fiber Optic,38.883224,-121.15918,1,68.6,0,9,Offer D,6096,0,0,1,0,15,2,111.0,362.55,0.0,1108.6,0,0,95658
6348,0,0,0,0,26,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),69.05,1815.65,0,49,30,37.51,5379,0,Nicolaus,0,0,Cable,38.788897999999996,-121.608624,0,69.05,0,0,None,751,0,0,0,0,26,1,0.0,975.26,0.0,1815.65,0,1,95659
6349,0,0,1,1,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.7,730.4,0,62,0,15.41,5636,0,North Highlands,0,0,NA,38.671295,-121.388251,1,19.7,2,5,None,32202,0,0,1,0,35,0,0.0,539.35,0.0,730.4,0,0,95660
6350,1,0,0,1,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.05,75.45,0,23,0,37.85,2948,0,Roseville,0,1,NA,38.736684999999994,-121.25198400000001,0,20.05,1,0,None,25173,0,0,0,0,3,0,0.0,113.55,0.0,75.45,1,0,95661
6351,1,0,1,1,50,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,103.7,5071.05,1,28,76,34.14,5897,1,Orangevale,0,1,Fiber Optic,38.689174,-121.21843500000001,1,107.848,0,1,Offer B,32040,1,1,1,1,50,3,3854.0,1707.0,36.61,5071.05,1,0,95662
6352,1,0,1,0,42,1,1,Fiber optic,1,0,0,1,Month-to-month,1,Electronic check,94.4,4014.6,0,52,11,41.16,2662,0,Penryn,1,1,Fiber Optic,38.859093,-121.182872,1,94.4,0,9,None,2048,0,0,1,1,42,0,442.0,1728.7199999999998,0.0,4014.6,0,0,95663
6353,1,0,1,0,10,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),54.95,568.85,0,34,9,21.85,3519,0,Pilot Hill,0,1,DSL,38.803731,-121.04379899999999,1,54.95,0,9,Offer D,1173,1,0,1,0,10,0,51.0,218.5,0.0,568.85,0,0,95664
6354,0,0,1,0,61,1,0,Fiber optic,1,1,0,1,One year,0,Bank transfer (automatic),93.7,5860.7,0,19,69,10.21,4300,0,Pine Grove,0,0,DSL,38.400264,-120.641274,1,93.7,0,0,None,4354,1,0,0,1,61,0,404.39,622.8100000000002,0.0,5860.7,1,1,95665
6355,0,0,0,0,68,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),110.25,7279.35,0,43,17,48.82,5502,0,Pioneer,0,0,Fiber Optic,38.546999,-120.27111399999998,0,110.25,0,0,None,5501,1,0,0,1,68,2,0.0,3319.76,0.0,7279.35,0,1,95666
6356,1,0,0,0,10,1,0,Fiber optic,1,0,1,1,One year,1,Electronic check,98.9,1064.95,0,37,26,46.33,4614,0,Placerville,1,1,DSL,38.733714,-120.79521299999999,0,98.9,0,0,Offer D,34146,0,1,0,1,10,1,0.0,463.3,0.0,1064.95,0,1,95667
6357,1,0,1,0,65,1,1,Fiber optic,1,1,0,0,One year,0,Electronic check,89.75,5769.6,1,39,18,49.33,6110,1,Pleasant Grove,1,1,Cable,38.833554,-121.498102,1,93.34,0,5,Offer B,901,0,2,1,0,65,4,0.0,3206.45,18.72,5769.6,0,1,95668
6358,0,0,1,1,72,1,0,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),80.45,5886.85,0,35,56,12.96,4480,0,Plymouth,1,0,Fiber Optic,38.489273,-120.89161399999999,1,80.45,3,3,None,2220,1,0,1,1,72,1,3297.0,933.12,0.0,5886.85,0,0,95669
6359,1,0,1,1,55,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Electronic check,79.4,4238.45,0,43,53,13.45,4162,0,Rancho Cordova,0,1,DSL,38.602723,-121.279913,1,79.4,3,9,None,49729,1,0,1,0,55,1,0.0,739.75,0.0,4238.45,0,1,95670
6360,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.3,20.3,1,44,0,26.37,3830,1,Rescue,0,0,NA,38.724321999999994,-120.99123700000001,0,20.3,0,0,Offer E,3815,0,0,0,0,1,2,0.0,26.37,0.0,20.3,0,0,95672
6361,0,0,0,0,7,1,0,DSL,0,0,0,1,Month-to-month,0,Bank transfer (automatic),62.8,418.3,0,42,21,8.29,4080,0,Rio Linda,1,0,DSL,38.688764,-121.457596,0,62.8,0,0,None,14010,1,0,0,1,7,0,88.0,58.03,0.0,418.3,0,0,95673
6362,0,0,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.9,136.05,0,50,25,41.08,2044,0,Rio Oso,0,0,Fiber Optic,38.954144,-121.48253600000001,0,74.9,0,0,None,947,0,0,0,0,2,1,34.0,82.16,0.0,136.05,0,0,95674
6363,0,0,0,0,9,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,74.85,708.2,0,28,73,13.05,5770,0,River Pines,0,0,DSL,38.545775,-120.743325,0,74.85,0,0,None,364,0,0,0,0,9,0,0.0,117.45,0.0,708.2,1,1,95675
6364,1,0,0,1,27,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.85,788.55,0,54,0,2.65,2682,0,Rocklin,0,1,NA,38.7904,-121.23697299999999,0,25.85,1,0,None,21510,0,0,0,0,27,1,0.0,71.55,0.0,788.55,0,0,95677
6365,1,1,1,0,7,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.95,700.85,1,65,3,34.66,2016,1,Roseville,1,1,Fiber Optic,38.759751,-121.288545,1,106.02799999999999,0,2,None,30614,0,0,1,1,7,0,0.0,242.62,0.0,700.85,0,1,95678
6366,0,0,1,0,64,1,0,DSL,0,1,0,1,Two year,1,Mailed check,68.3,4378.8,0,57,25,23.29,5425,0,Sheridan,1,0,Cable,38.984756,-121.345074,1,68.3,0,9,None,1219,1,0,1,1,64,1,1095.0,1490.56,0.0,4378.8,0,0,95681
6367,1,0,0,0,70,0,No phone service,DSL,1,0,0,1,Two year,0,Bank transfer (automatic),48.4,3442.8,0,23,26,0.0,4483,0,Shingle Springs,1,1,Fiber Optic,38.598936,-120.96309199999999,0,48.4,0,0,None,24738,1,0,0,1,70,0,0.0,0.0,0.0,3442.8,1,1,95682
6368,1,1,0,0,2,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.0,181.7,1,65,24,20.99,5569,1,Sloughhouse,0,1,DSL,38.470423,-121.114897,0,97.76,0,0,Offer E,4731,0,0,0,1,2,2,4.36,41.98,0.0,181.7,0,1,95683
6369,1,1,0,0,67,1,0,Fiber optic,1,1,1,1,Two year,1,Electronic check,105.05,7171.7,0,65,11,34.23,4143,0,Somerset,0,1,Fiber Optic,38.606703,-120.58665900000001,0,105.05,0,0,None,2958,1,0,0,1,67,1,789.0,2293.41,0.0,7171.7,0,0,95684
6370,0,0,0,0,45,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),89.3,4016.85,1,41,26,14.12,4880,1,Sutter Creek,0,0,Cable,38.432145,-120.77068999999999,0,92.87200000000001,0,0,Offer B,4610,0,0,0,0,45,8,1044.0,635.4,44.63,4016.85,0,0,95685
6371,0,0,0,0,24,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.15,553,0,19,0,26.64,3904,0,Thornton,0,0,NA,38.157794,-121.520223,0,25.15,0,0,None,1472,0,0,0,0,24,1,0.0,639.36,0.0,553.0,1,0,95686
6372,1,0,1,1,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.5,96.85,0,62,0,3.57,5390,0,Vacaville,0,1,NA,38.333133000000004,-121.920151,1,19.5,2,8,None,63157,0,1,1,0,4,1,0.0,14.28,0.0,96.85,0,0,95687
6373,1,0,1,1,44,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),92.95,4122.9,0,46,25,26.25,5635,0,Vacaville,1,1,Fiber Optic,38.419088,-122.02456799999999,1,92.95,1,2,None,32564,0,0,1,1,44,0,1031.0,1155.0,0.0,4122.9,0,0,95688
6374,0,0,1,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.7,1482.3,0,64,0,6.9,4528,0,Volcano,0,0,NA,38.481902000000005,-120.603668,1,20.7,3,9,None,1273,0,0,1,0,72,2,0.0,496.8,0.0,1482.3,0,0,95689
6375,0,0,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),74.3,74.3,1,31,9,39.66,5996,1,Walnut Grove,0,0,Cable,38.240419,-121.587535,0,77.27199999999999,0,0,Offer E,2344,0,0,0,0,1,0,0.0,39.66,0.0,74.3,0,1,95690
6376,1,0,0,0,66,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.35,1240.8,0,58,0,21.23,5637,0,West Sacramento,0,1,NA,38.627951,-121.59328700000002,0,19.35,0,0,None,19050,0,0,0,0,66,1,0.0,1401.18,0.0,1240.8,0,0,95691
6377,1,0,0,0,1,0,No phone service,DSL,0,1,0,1,Month-to-month,1,Mailed check,44.65,44.65,1,49,21,0.0,3704,1,Wheatland,0,1,Cable,39.043387,-121.40983700000001,0,46.43600000000001,0,0,Offer E,3600,1,1,0,1,1,4,0.0,0.0,0.0,44.65,0,1,95692
6378,1,0,1,1,13,1,0,Fiber optic,1,0,0,1,Month-to-month,0,Electronic check,84.05,1095.3,1,40,23,29.92,4745,1,Wilton,0,1,Fiber Optic,38.392559000000006,-121.22509299999999,1,87.412,0,5,Offer D,5889,0,0,1,1,13,2,25.19,388.96,23.97,1095.3,0,1,95693
6379,1,0,0,0,10,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),80.7,788.8,1,54,3,17.07,3492,1,Winters,0,1,Fiber Optic,38.578604,-122.024579,0,83.92800000000003,0,0,Offer D,8406,0,0,0,0,10,2,0.0,170.7,38.42,788.8,0,1,95694
6380,1,1,1,0,65,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,104.35,6578.55,0,76,7,8.59,4073,0,Woodland,1,1,Fiber Optic,38.71967,-121.862416,1,104.35,0,9,Offer B,38547,0,0,1,0,65,0,0.0,558.35,0.0,6578.55,0,1,95695
6381,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.55,19.55,0,42,0,30.63,5272,0,Alta,0,1,NA,39.218096,-120.79153000000001,0,19.55,3,0,None,751,0,0,0,0,1,3,0.0,30.63,0.0,19.55,0,0,95701
6382,1,0,1,1,38,1,0,DSL,1,1,1,0,One year,0,Electronic check,74.05,2802.3,0,59,76,31.45,5975,0,Applegate,1,1,Fiber Optic,38.983388,-120.98881399999999,1,74.05,3,4,None,1526,1,0,1,0,38,1,0.0,1195.1,0.0,2802.3,0,1,95703
6383,1,0,0,1,23,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,40.1,857.75,0,36,26,0.0,2327,0,Camino,1,1,DSL,38.748315999999996,-120.67551200000001,0,40.1,3,0,None,4829,1,0,0,0,23,0,223.0,0.0,0.0,857.75,0,0,95709
6384,0,0,1,0,10,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,184.4,0,23,0,14.04,3509,0,Colfax,0,0,NA,39.084645,-120.89401399999998,1,20.1,0,4,None,8525,0,0,1,0,10,1,0.0,140.39999999999998,0.0,184.4,1,0,95713
6385,1,0,0,1,4,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.7,364.55,1,28,94,26.16,2777,1,Dutch Flat,0,1,Cable,39.197215,-120.83679,0,105.76799999999999,0,0,Offer E,350,0,0,0,1,4,3,343.0,104.64,1.48,364.55,1,0,95714
6386,1,0,1,1,72,1,1,DSL,1,0,1,1,Two year,1,Credit card (automatic),83.55,6093.3,0,25,27,21.21,5940,0,Emigrant Gap,1,1,Cable,39.23754,-120.720196,1,83.55,2,4,None,185,1,1,1,1,72,1,0.0,1527.12,0.0,6093.3,1,1,95715
6387,0,0,1,0,35,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,56.85,1861.1,0,20,69,20.79,3102,0,Gold Run,0,0,Fiber Optic,39.170376,-120.838404,1,56.85,0,7,None,407,1,0,1,0,35,2,1284.0,727.65,0.0,1861.1,1,0,95717
6388,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,20.4,1,31,0,22.12,3663,1,Kyburz,0,0,NA,38.766036,-120.209673,0,20.4,0,0,Offer E,183,0,0,0,0,1,1,0.0,22.12,0.0,20.4,0,0,95720
6389,0,0,1,1,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.55,1079.65,0,52,0,43.52,4125,0,Echo Lake,0,0,NA,38.851842,-120.076204,1,19.55,2,4,None,69,0,0,1,0,58,1,0.0,2524.1600000000008,0.0,1079.65,0,0,95721
6390,1,0,1,1,70,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,106.15,7475.1,0,37,28,3.67,4649,0,Meadow Vista,1,1,Fiber Optic,39.003358,-121.022539,1,106.15,3,7,None,3747,1,0,1,1,70,1,2093.0,256.9,0.0,7475.1,0,0,95722
6391,1,0,1,1,38,1,1,DSL,0,1,1,1,One year,0,Credit card (automatic),78.95,2862.55,0,56,30,13.67,2125,0,Pollock Pines,1,1,Fiber Optic,38.733908,-120.45341599999999,1,78.95,3,2,None,8577,0,1,1,1,38,1,859.0,519.46,0.0,2862.55,0,0,95726
6392,0,0,1,1,60,0,No phone service,DSL,0,1,1,1,Month-to-month,1,Electronic check,49.75,3069.45,0,39,51,0.0,6307,0,Soda Springs,0,0,Fiber Optic,39.279068,-120.414275,1,49.75,3,2,None,88,0,0,1,1,60,1,1565.0,0.0,0.0,3069.45,0,0,95728
6393,1,0,0,0,26,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Credit card (automatic),92.4,2349.8,0,34,8,37.59,5461,0,Twin Bridges,0,1,Cable,38.805481,-120.13287,0,92.4,0,0,None,25,0,0,0,0,26,2,0.0,977.34,0.0,2349.8,0,1,95735
6394,0,0,0,0,8,1,0,DSL,1,1,0,0,One year,0,Bank transfer (automatic),58.2,469.25,0,60,28,17.52,3325,0,Weimar,0,0,Cable,39.00978,-120.978273,0,58.2,0,0,None,31,1,0,0,0,8,2,0.0,140.16,0.0,469.25,0,1,95736
6395,1,0,1,1,41,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,102.6,4213.35,1,36,11,45.03,2098,1,Rancho Cordova,1,1,Cable,38.591134000000004,-121.161585,1,106.704,0,1,Offer B,299,1,2,1,1,41,4,463.0,1846.23,2.93,4213.35,0,0,95742
6396,0,1,1,0,36,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),91.95,3301.05,0,74,16,11.32,3273,0,Granite Bay,0,0,DSL,38.749466,-121.184196,1,91.95,0,0,Offer C,20675,0,0,0,0,36,0,0.0,407.52,17.76,3301.05,0,1,95746
6397,1,1,0,0,54,1,0,DSL,0,0,0,1,One year,0,Bank transfer (automatic),65.25,3529.95,0,79,6,5.14,6161,0,Roseville,1,1,Fiber Optic,38.784329,-121.373245,0,65.25,0,0,Offer B,25418,1,0,0,0,54,2,212.0,277.56,33.07,3529.95,0,0,95747
6398,1,0,1,1,71,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),106.0,7723.7,1,60,13,47.34,4072,1,Elk Grove,1,1,Cable,38.353629999999995,-121.44195,1,110.24,0,3,Offer A,47065,0,0,1,1,71,4,1004.0,3361.140000000001,0.0,7723.7,0,0,95758
6399,0,0,0,0,55,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.1,4144.9,0,50,26,8.93,5832,0,El Dorado Hills,0,0,Fiber Optic,38.684437,-121.05563400000001,0,73.1,0,0,None,22028,0,0,0,0,55,2,1078.0,491.15,0.0,4144.9,0,0,95762
6400,0,0,0,0,72,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),59.75,4265,0,40,23,12.63,4515,0,Rocklin,0,0,Fiber Optic,38.823278,-121.281856,0,59.75,0,0,None,15494,0,0,0,0,72,0,0.0,909.36,0.0,4265.0,0,1,95765
6401,0,0,0,1,3,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,55.1,154.65,1,43,18,26.04,4412,1,Woodland,0,0,Cable,38.694081,-121.69443100000001,0,57.303999999999995,2,0,Offer E,15022,1,0,0,0,3,4,28.0,78.12,0.0,154.65,0,0,95776
6402,0,0,1,1,54,1,1,DSL,0,1,0,0,Two year,1,Bank transfer (automatic),59.8,3246.45,0,61,21,23.02,5898,0,Sacramento,1,0,DSL,38.584505,-121.491956,1,59.8,3,9,None,16599,0,0,1,0,54,0,0.0,1243.08,0.0,3246.45,0,1,95814
6403,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),116.6,8337.45,0,26,52,21.29,5227,0,Sacramento,1,1,Fiber Optic,38.608405,-121.449942,1,116.6,1,7,None,25355,1,0,1,1,72,0,0.0,1532.88,26.7,8337.45,1,1,95815
6404,1,0,0,0,52,1,1,Fiber optic,1,0,1,1,Two year,1,Electronic check,109.3,5731.4,0,54,30,20.8,5624,0,Sacramento,1,1,Fiber Optic,38.574856,-121.46503999999999,0,109.3,0,0,None,16164,1,0,0,1,52,0,0.0,1081.6,3.85,5731.4,0,1,95816
6405,0,1,0,0,60,1,1,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),101.4,6176.6,0,74,11,48.92,4483,0,Sacramento,0,0,Cable,38.550722,-121.457314,0,101.4,0,0,Offer B,14966,0,0,0,0,60,0,679.0,2935.2000000000007,0.0,6176.6,0,0,95817
6406,0,0,0,0,39,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),50.65,1905.4,0,56,6,0.0,5433,0,Sacramento,1,0,DSL,38.556306,-121.49581699999999,0,50.65,0,0,None,21313,0,0,0,1,39,0,11.43,0.0,3.51,1905.4,0,1,95818
6407,0,0,0,0,15,1,0,DSL,0,0,1,0,One year,0,Mailed check,56.15,931.9,0,28,52,6.56,5473,0,Sacramento,0,0,DSL,38.567594,-121.43750700000001,0,56.15,0,0,None,15975,0,0,0,0,15,2,485.0,98.4,35.23,931.9,1,0,95819
6408,1,0,0,0,69,1,1,Fiber optic,0,0,1,1,Two year,1,Bank transfer (automatic),106.5,7348.8,1,58,12,26.88,4859,1,Sacramento,1,1,Cable,38.53508,-121.444144,0,110.76,0,0,Offer A,37031,1,0,0,1,69,1,882.0,1854.72,0.0,7348.8,0,0,95820
6409,1,0,1,1,43,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.2,776.25,0,39,0,14.97,5594,0,Sacramento,0,1,NA,38.625096,-121.38365800000001,1,19.2,1,10,None,35426,0,0,1,0,43,2,0.0,643.71,9.48,776.25,0,0,95821
6410,0,1,0,0,63,1,1,DSL,1,1,1,0,One year,0,Bank transfer (automatic),83.0,5243.05,0,71,18,15.62,5428,0,Sacramento,1,0,DSL,38.512569,-121.49518400000001,0,83.0,0,0,Offer B,44683,1,0,0,0,63,2,944.0,984.06,0.0,5243.05,0,0,95822
6411,1,1,1,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.1,141.65,0,70,24,34.99,5592,0,Sacramento,0,1,DSL,38.475465,-121.443625,1,70.1,0,9,Offer E,72199,0,0,1,0,2,3,34.0,69.98,0.0,141.65,0,0,95823
6412,0,0,1,1,72,1,0,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),108.3,7679.65,0,51,25,41.55,4183,0,Sacramento,1,0,Fiber Optic,38.517295000000004,-121.439819,1,108.3,2,1,None,30580,1,0,1,1,72,1,1920.0,2991.6,36.13,7679.65,0,0,95824
6413,0,0,1,1,32,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),91.05,2954.5,1,51,10,46.92,3590,1,Sacramento,1,0,Cable,38.590035,-121.41245500000001,1,94.692,0,1,None,30715,0,1,1,1,32,5,295.0,1501.44,0.0,2954.5,0,0,95825
6414,1,0,1,1,40,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.25,1006.9,0,43,0,27.95,3217,0,Sacramento,0,1,NA,38.542532,-121.378826,1,25.25,1,9,None,38818,0,0,1,0,40,0,0.0,1118.0,44.51,1006.9,0,0,95826
6415,0,0,1,0,58,0,No phone service,DSL,1,1,1,0,One year,1,Electronic check,45.35,2540.1,0,55,29,0.0,5137,0,Sacramento,0,0,Fiber Optic,38.549184999999994,-121.32838600000001,1,45.35,0,7,None,19611,0,0,1,0,58,0,737.0,0.0,4.08,2540.1,0,0,95827
6416,1,0,0,0,67,0,No phone service,DSL,1,0,1,0,Two year,0,Electronic check,43.9,3097.2,0,44,17,0.0,6344,0,Sacramento,0,1,Fiber Optic,38.486938,-121.39580500000001,0,43.9,0,0,None,54880,1,0,0,0,67,0,527.0,0.0,34.45,3097.2,0,0,95828
6417,0,1,1,0,51,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Electronic check,77.5,3807.35,1,69,10,17.87,5748,1,Sacramento,0,0,Cable,38.486502,-121.334051,1,80.60000000000002,0,1,None,11396,0,0,1,0,51,7,381.0,911.37,0.0,3807.35,0,0,95829
6418,1,0,1,0,31,1,1,DSL,0,0,1,1,One year,1,Mailed check,79.3,2484,0,47,6,3.12,5238,0,Sacramento,1,1,DSL,38.490508,-121.284171,1,79.3,0,1,None,592,1,0,1,1,31,0,14.9,96.72,0.0,2484.0,0,1,95830
6419,1,1,1,0,69,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),84.9,5785.65,0,77,14,14.76,4503,0,Sacramento,0,1,DSL,38.494832,-121.52944699999999,1,84.9,0,7,None,42832,0,0,1,0,69,1,810.0,1018.44,0.0,5785.65,0,0,95831
6420,1,0,1,0,32,1,1,Fiber optic,0,0,0,0,One year,1,Electronic check,79.25,2619.15,0,64,18,43.11,2735,0,Sacramento,0,1,Fiber Optic,38.445939,-121.49685500000001,1,79.25,0,4,None,9063,1,0,1,0,32,0,471.0,1379.52,16.96,2619.15,0,0,95832
6421,0,0,0,0,21,1,0,DSL,1,1,1,0,Two year,0,Credit card (automatic),71.05,1524.85,0,23,71,17.35,5138,0,Sacramento,0,0,DSL,38.619049,-121.517552,0,71.05,0,0,None,31422,1,0,0,0,21,0,0.0,364.35,16.91,1524.85,1,1,95833
6422,1,0,0,0,52,1,0,DSL,1,0,0,0,One year,0,Electronic check,53.75,2790.65,0,42,3,47.9,5957,0,Sacramento,1,1,Cable,38.646209000000006,-121.52446,0,53.75,0,0,None,8403,0,0,0,0,52,1,0.0,2490.8,43.12,2790.65,0,1,95834
6423,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),24.25,1784.5,0,42,0,47.6,5897,0,Sacramento,0,0,NA,38.685069,-121.543709,1,24.25,3,8,None,854,0,0,1,0,72,1,0.0,3427.2000000000007,49.76,1784.5,0,0,95835
6424,0,0,1,0,72,0,No phone service,DSL,0,1,1,1,Two year,1,Electronic check,54.2,3937.45,1,51,16,0.0,4481,1,Sacramento,1,0,Cable,38.691607,-121.60228400000001,1,56.368,0,1,Offer A,264,0,0,1,1,72,2,630.0,0.0,0.0,3937.45,0,0,95837
6425,1,0,1,1,52,0,No phone service,DSL,1,0,0,1,One year,0,Bank transfer (automatic),44.25,2276.1,0,48,19,0.0,6340,0,Sacramento,1,1,Fiber Optic,38.646096,-121.44243300000001,1,44.25,2,9,None,34894,0,0,1,1,52,1,432.0,0.0,23.5,2276.1,0,0,95838
6426,0,0,0,0,41,1,0,DSL,0,0,0,0,One year,0,Bank transfer (automatic),50.05,2029.05,0,62,12,12.42,2157,0,Sacramento,0,0,Cable,38.660441999999996,-121.346321,0,50.05,0,0,None,20993,1,0,0,0,41,3,243.0,509.22,0.0,2029.05,0,0,95841
6427,1,0,0,0,41,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.15,802.35,0,46,0,36.76,4982,0,Sacramento,0,1,NA,38.687367,-121.34848000000001,0,20.15,0,0,None,31373,0,0,0,0,41,0,0.0,1507.16,29.95,802.35,0,0,95842
6428,0,0,0,0,6,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.25,418.4,1,50,6,39.36,5816,1,Antelope,0,0,DSL,38.715498,-121.36341100000001,0,72.02,0,0,None,36432,0,0,0,0,6,3,0.0,236.16,0.0,418.4,0,1,95843
6429,1,0,1,1,67,1,1,DSL,1,1,0,0,One year,1,Credit card (automatic),69.35,4653.25,0,39,24,36.21,5589,0,Sacramento,1,1,Fiber Optic,38.585826000000004,-121.376263,1,69.35,1,6,None,23362,1,1,1,0,67,2,111.68,2426.07,9.99,4653.25,0,1,95864
6430,0,0,1,1,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.35,275.9,0,40,0,12.82,4146,0,Marysville,0,0,NA,39.19514,-121.503883,1,19.35,3,10,None,38091,0,0,1,0,16,1,0.0,205.12,33.24,275.9,0,0,95901
6431,1,0,0,0,17,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.15,343.45,0,35,0,27.66,2717,0,Beale Afb,0,1,NA,39.125310999999996,-121.392283,0,19.15,0,0,None,5654,0,0,0,0,17,2,0.0,470.22,28.63,343.45,0,0,95903
6432,1,0,1,0,35,1,0,DSL,1,1,0,0,Month-to-month,0,Mailed check,61.0,2130.45,0,27,30,25.32,4355,0,Alleghany,1,1,DSL,39.467828000000004,-120.84138600000001,1,61.0,0,4,None,118,0,0,1,0,35,2,0.0,886.2,10.7,2130.45,1,1,95910
6433,0,0,1,1,58,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.5,1191.4,0,52,0,25.86,6186,0,Arbuckle,0,0,NA,38.982372999999995,-122.047751,1,20.5,2,10,None,4796,0,0,1,0,58,1,0.0,1499.88,36.92,1191.4,0,0,95912
6434,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,50.5,50.5,1,35,31,39.58,2077,1,Bangor,1,1,Fiber Optic,39.396584999999995,-121.38028999999999,0,52.52,0,0,None,626,0,0,0,0,1,5,0.0,39.58,0.0,50.5,0,1,95914
6435,1,0,1,1,52,0,No phone service,DSL,0,1,1,0,Two year,0,Mailed check,50.2,2554,0,35,17,0.0,5396,0,Berry Creek,1,1,Cable,39.657228,-121.37778,1,50.2,2,1,None,1279,1,0,1,0,52,0,434.0,0.0,27.01,2554.0,0,0,95916
6436,0,0,0,0,70,1,0,DSL,1,0,1,1,Two year,0,Bank transfer (automatic),79.6,5589.45,0,60,28,47.72,5474,0,Biggs,1,0,Cable,39.457388,-121.818201,0,79.6,0,0,None,3169,1,0,0,1,70,2,1565.0,3340.4,42.34,5589.45,0,0,95917
6437,0,0,1,1,19,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),24.9,467.7,0,20,0,31.58,5396,0,Browns Valley,0,0,NA,39.292334000000004,-121.32059699999999,1,24.9,1,1,None,1477,0,1,1,0,19,1,0.0,600.02,0.0,467.7,1,0,95918
6438,1,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.4,74.4,1,68,13,11.08,3429,1,Brownsville,0,1,Fiber Optic,39.440687,-121.26358300000001,0,77.376,0,0,Offer E,1237,0,0,0,0,1,1,0.0,11.08,0.0,74.4,0,0,95919
6439,0,0,1,1,35,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,106.9,3756.45,0,33,56,26.09,5447,0,Butte City,1,0,Cable,39.449794,-121.93637199999999,1,106.9,3,1,None,303,1,0,1,1,35,0,0.0,913.15,34.47,3756.45,0,1,95920
6440,0,0,0,0,32,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.35,3334.9,0,33,28,41.53,4341,0,Camptonville,1,0,DSL,39.432127,-121.09928700000002,0,101.35,0,0,None,632,0,0,0,1,32,0,934.0,1328.96,0.0,3334.9,0,0,95922
6441,0,0,1,1,17,1,0,DSL,1,0,0,0,Month-to-month,1,Credit card (automatic),55.35,920.5,0,25,69,20.23,5465,0,Canyon Dam,0,0,DSL,40.171312,-121.120605,1,55.35,3,1,None,86,1,0,1,0,17,1,0.0,343.91,0.0,920.5,1,1,95923
6442,0,0,1,1,67,1,0,DSL,0,1,0,0,One year,0,Credit card (automatic),50.55,3431.75,0,44,28,46.9,5122,0,Challenge,0,0,Fiber Optic,39.461768,-121.195825,1,50.55,3,1,Offer A,262,0,0,1,0,67,2,961.0,3142.3,0.0,3431.75,0,0,95925
6443,0,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.5,150.35,0,56,0,43.83,4883,0,Chico,0,0,NA,39.745712,-121.84333000000001,0,19.5,0,0,None,35808,0,0,0,0,9,3,0.0,394.47,0.0,150.35,0,0,95926
6444,1,0,0,1,31,1,1,DSL,0,1,1,1,One year,1,Mailed check,79.45,2587.7,1,37,3,6.71,2872,1,Chico,0,1,DSL,39.681488,-121.83721000000001,0,82.62799999999999,0,0,None,32848,1,1,0,1,31,2,78.0,208.01,0.0,2587.7,0,0,95928
6445,1,0,0,0,4,1,1,Fiber optic,1,0,1,0,Month-to-month,0,Electronic check,90.65,367.95,0,43,18,31.57,3559,0,Clipper Mills,0,1,Cable,39.562239,-121.14836000000001,0,90.65,0,0,Offer E,282,0,0,0,0,4,0,66.0,126.28,0.0,367.95,0,0,95930
6446,1,1,1,1,58,1,1,Fiber optic,1,1,0,0,One year,1,Bank transfer (automatic),89.85,5125.75,0,71,10,18.43,5035,0,Colusa,0,1,Fiber Optic,39.273096,-122.05076299999999,1,89.85,1,1,Offer B,7503,1,0,1,0,58,0,0.0,1068.94,0.0,5125.75,0,1,95932
6447,1,0,0,0,60,1,0,DSL,1,0,1,1,One year,0,Mailed check,79.0,4801.1,0,62,3,35.13,4807,0,Crescent Mills,1,1,Cable,40.080342,-120.95780500000001,0,79.0,0,0,None,178,1,0,0,1,60,0,0.0,2107.8,0.0,4801.1,0,1,95934
6448,1,0,0,0,58,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,104.65,6219.6,1,34,28,41.14,5411,1,Dobbins,1,1,Fiber Optic,39.381174,-121.21191,0,108.836,0,0,Offer B,614,1,1,0,1,58,2,1741.0,2386.12,0.0,6219.6,0,0,95935
6449,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.55,19.55,0,35,0,17.94,3718,0,Downieville,0,1,NA,39.578792,-120.780786,0,19.55,0,0,Offer E,404,0,0,0,0,1,1,0.0,17.94,0.0,19.55,0,0,95936
6450,0,0,1,1,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.9,550.1,0,36,0,2.4,4870,0,Dunnigan,0,0,NA,38.931425,-121.946081,1,19.9,3,1,None,19,0,0,1,0,27,0,0.0,64.8,0.0,550.1,0,0,95937
6451,1,1,1,1,66,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,116.25,7862.25,0,77,10,3.27,4578,0,Durham,1,1,Fiber Optic,39.607831,-121.77795900000001,1,116.25,2,0,None,3524,1,0,0,0,66,3,0.0,215.82,0.0,7862.25,0,1,95938
6452,1,0,0,0,15,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Bank transfer (automatic),87.75,1242.2,0,20,59,13.8,5415,0,Elk Creek,0,1,Fiber Optic,39.53222,-122.594879,0,87.75,0,0,None,587,0,0,0,0,15,1,733.0,207.0,0.0,1242.2,1,0,95939
6453,1,1,1,0,47,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.05,4871.05,1,68,21,8.97,5166,1,Forbestown,1,1,DSL,39.531028000000006,-121.24807,1,104.052,0,1,None,452,0,0,1,0,47,2,1023.0,421.59,0.0,4871.05,0,0,95941
6454,0,0,0,0,41,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),81.3,3190.65,0,32,19,7.83,2299,0,Forest Ranch,0,0,Fiber Optic,40.077028000000006,-121.49416799999999,0,81.3,0,0,None,1351,0,1,0,0,41,1,0.0,321.0300000000001,0.0,3190.65,0,1,95942
6455,1,0,1,0,59,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,44.3,2666.75,0,21,53,0.0,5905,0,Glenn,0,1,DSL,39.597975,-122.032248,1,44.3,0,1,Offer B,1454,0,0,1,1,59,0,0.0,0.0,0.0,2666.75,1,1,95943
6456,0,0,0,1,50,1,0,Fiber optic,0,0,0,0,Two year,0,Credit card (automatic),70.35,3533.6,0,45,20,36.11,5521,0,Goodyears Bar,0,0,DSL,39.564113,-120.86883600000002,0,70.35,2,0,Offer B,76,0,0,0,0,50,2,0.0,1805.5,0.0,3533.6,0,1,95944
6457,1,0,1,1,17,0,No phone service,DSL,1,0,1,0,One year,0,Credit card (automatic),44.45,792.15,0,20,52,0.0,3522,0,Grass Valley,1,1,Cable,39.194539,-120.98806599999999,1,44.45,2,1,None,23990,0,0,1,0,17,3,0.0,0.0,0.0,792.15,1,1,95945
6458,1,0,1,1,6,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.15,295.65,0,48,51,34.7,4076,0,Penn Valley,0,1,DSL,39.203817,-121.19583999999999,1,49.15,3,1,Offer E,9752,0,0,1,0,6,1,0.0,208.2,0.0,295.65,0,1,95946
6459,1,1,1,0,51,0,No phone service,DSL,0,1,0,0,Month-to-month,1,Credit card (automatic),29.45,1459.35,0,71,21,0.0,6285,0,Greenville,0,1,Fiber Optic,40.160385999999995,-120.83542800000001,1,29.45,0,1,Offer B,2064,0,0,1,0,51,0,306.0,0.0,0.0,1459.35,0,0,95947
6460,1,0,0,0,44,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,100.55,4398.15,1,41,25,42.92,3486,1,Gridley,0,1,Cable,39.346897999999996,-121.75953700000001,0,104.572,0,0,None,9763,1,2,0,1,44,4,1100.0,1888.48,0.0,4398.15,0,0,95948
6461,1,0,1,0,49,1,0,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),85.3,4297.95,0,44,23,14.21,4696,0,Grass Valley,0,1,Fiber Optic,39.099204,-121.13796200000002,1,85.3,0,1,Offer B,17922,0,0,1,0,49,2,989.0,696.2900000000002,0.0,4297.95,0,0,95949
6462,1,0,0,0,2,1,0,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,95.65,167.3,1,34,30,16.76,5332,1,Grimes,0,1,Cable,39.033058000000004,-121.89571799999999,0,99.476,0,0,None,531,0,0,0,1,2,3,50.0,33.52,0.0,167.3,0,0,95950
6463,1,0,1,0,59,1,1,DSL,1,0,0,1,One year,1,Mailed check,69.1,4096.9,0,30,53,20.5,4765,0,Hamilton City,0,1,Fiber Optic,39.732766999999996,-122.042298,1,69.1,0,1,Offer B,1931,1,0,1,1,59,0,2171.0,1209.5,0.0,4096.9,0,0,95951
6464,1,1,0,0,50,1,1,DSL,1,1,1,0,Month-to-month,1,Bank transfer (automatic),70.35,3454.6,0,69,23,25.23,5596,0,Live Oak,0,1,Fiber Optic,39.258746,-121.77696999999999,0,70.35,0,0,Offer B,8695,0,0,0,0,50,2,795.0,1261.5,0.0,3454.6,0,0,95953
6465,0,0,1,1,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.6,1286,0,45,0,2.47,6325,0,Magalia,0,0,NA,39.933852,-121.58437099999999,1,20.6,2,1,Offer B,11168,0,0,1,0,59,0,0.0,145.73000000000005,0.0,1286.0,0,0,95954
6466,1,0,0,0,18,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,74.15,1387,0,63,20,4.38,2643,0,Maxwell,0,1,Fiber Optic,39.281194,-122.226568,0,74.15,0,0,None,1146,0,0,0,0,18,2,277.0,78.84,0.0,1387.0,0,0,95955
6467,1,0,0,0,10,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,75.05,786.3,0,22,26,17.98,3399,0,Meadow Valley,0,1,Cable,39.937017,-121.058043,0,75.05,0,0,None,301,0,0,0,0,10,1,0.0,179.8,0.0,786.3,1,1,95956
6468,1,0,1,0,14,1,0,DSL,0,0,0,0,One year,0,Electronic check,44.6,641.25,0,57,19,44.95,4612,0,Meridian,0,1,DSL,39.068071,-121.83263799999999,1,44.6,0,1,Offer D,776,0,0,1,0,14,0,122.0,629.3000000000002,0.0,641.25,0,0,95957
6469,1,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),21.45,705.45,0,47,0,17.2,3967,0,Nevada City,0,1,NA,39.333737,-120.858667,0,21.45,0,0,None,17269,0,0,0,0,35,1,0.0,602.0,0.0,705.45,0,0,95959
6470,1,0,1,1,8,1,0,DSL,0,0,0,0,One year,1,Mailed check,43.45,345.5,0,48,24,6.78,4184,0,North San Juan,0,1,Fiber Optic,39.423046,-120.984472,1,43.45,2,1,Offer E,565,0,0,1,0,8,1,0.0,54.24,0.0,345.5,0,1,95960
6471,1,0,1,1,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.05,345.9,0,56,0,28.06,4458,0,Olivehurst,0,1,NA,39.082568,-121.55325,1,20.05,3,1,Offer D,6439,0,0,1,0,18,1,0.0,505.08,0.0,345.9,0,0,95961
6472,0,0,1,1,60,1,1,Fiber optic,1,1,1,0,One year,0,Bank transfer (automatic),94.15,5811.8,0,35,76,48.04,6399,0,Oregon House,0,0,Cable,39.342587,-121.24983300000001,1,94.15,3,1,Offer B,1519,0,0,1,0,60,0,441.7,2882.4,0.0,5811.8,0,1,95962
6473,0,0,0,0,1,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,94.4,94.4,1,49,7,18.34,5764,1,Orland,1,0,Cable,39.748037,-122.30216899999999,0,98.17600000000002,0,0,None,13706,0,0,0,1,1,2,0.0,18.34,0.0,94.4,0,0,95963
6474,0,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.55,124.45,0,61,0,7.35,5980,0,Oroville,0,0,NA,39.624561,-121.552866,0,19.55,0,0,Offer E,17782,0,0,0,0,6,2,0.0,44.1,0.0,124.45,0,0,95965
6475,0,0,0,1,19,1,1,DSL,1,1,1,0,Month-to-month,1,Mailed check,75.9,1375.6,0,49,57,8.02,4198,0,Oroville,0,0,Cable,39.473896,-121.415927,0,75.9,3,0,Offer D,28382,1,0,0,0,19,1,784.0,152.38,0.0,1375.6,0,0,95966
6476,1,0,1,1,53,1,1,DSL,1,1,0,0,One year,0,Bank transfer (automatic),64.15,3491.55,0,35,15,37.57,5570,0,Palermo,0,1,Fiber Optic,39.435756,-121.552071,1,64.15,2,1,Offer B,1254,1,0,1,0,53,0,524.0,1991.21,0.0,3491.55,0,0,95968
6477,1,1,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,1,Bank transfer (automatic),109.55,7920.7,0,67,4,17.71,4086,0,Paradise,1,1,Fiber Optic,39.69676,-121.644379,1,109.55,0,1,None,28318,0,0,1,1,72,0,0.0,1275.12,0.0,7920.7,0,1,95969
6478,0,0,1,0,60,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),110.8,6640.7,0,34,14,30.23,5942,0,Princeton,1,0,Fiber Optic,39.424957,-122.03930700000001,1,110.8,0,1,Offer B,495,1,0,1,1,60,0,930.0,1813.8,9.79,6640.7,0,0,95970
6479,0,0,0,0,1,1,0,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),55.0,55,1,47,29,32.74,3809,1,Quincy,0,0,Cable,39.971228,-121.04116599999999,0,57.2,0,0,None,6189,0,0,0,0,1,8,0.0,32.74,0.0,55.0,0,0,95971
6480,0,0,0,1,13,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,53.45,718.1,0,40,27,25.33,4335,0,Chico,1,0,Fiber Optic,39.903271999999994,-121.843567,0,53.45,1,0,Offer D,26971,1,1,0,0,13,1,0.0,329.29,26.37,718.1,0,1,95973
6481,0,0,1,1,5,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Credit card (automatic),69.95,320.4,0,47,16,1.38,3850,0,Richvale,0,0,DSL,39.495768,-121.747472,1,69.95,2,1,None,74,0,0,1,0,5,0,0.0,6.9,0.0,320.4,0,1,95974
6482,1,0,0,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,101.45,101.45,1,32,8,10.38,4390,1,Rough And Ready,1,1,Cable,39.225634,-121.15616299999999,0,105.508,0,0,None,1601,0,0,0,1,1,3,0.0,10.38,0.0,101.45,0,1,95975
6483,1,0,1,1,13,1,0,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,97.0,1334.45,0,60,19,44.05,5282,0,Smartville,1,1,DSL,39.176595,-121.291692,1,97.0,1,1,Offer D,963,0,0,1,1,13,0,0.0,572.65,0.0,1334.45,0,1,95977
6484,1,0,0,0,37,1,1,DSL,1,1,1,1,One year,1,Bank transfer (automatic),90.6,3358.65,0,42,6,44.52,2546,0,Stirling City,1,1,Fiber Optic,39.904002,-121.527823,0,90.6,0,0,None,28,1,0,0,1,37,2,0.0,1647.24,8.96,3358.65,0,1,95978
6485,1,0,1,0,64,1,0,Fiber optic,1,0,0,0,Month-to-month,1,Mailed check,73.55,4764,0,40,22,48.41,5018,0,Stonyford,0,1,Fiber Optic,39.288127,-122.41584099999999,1,73.55,0,0,Offer B,844,0,0,0,0,64,1,0.0,3098.24,21.9,4764.0,0,1,95979
6486,0,0,1,0,5,1,1,DSL,0,0,1,0,Month-to-month,0,Bank transfer (automatic),67.95,350.3,1,39,4,14.9,3889,1,Strawberry Valley,1,0,Cable,39.584579999999995,-121.09325600000001,1,70.668,0,1,None,101,1,0,1,0,5,1,0.0,74.5,0.0,350.3,0,1,95981
6487,0,0,1,0,61,1,1,Fiber optic,0,1,0,1,Two year,1,Bank transfer (automatic),94.35,5703,0,55,13,25.14,4676,0,Sutter,0,0,DSL,39.172777,-121.80584499999999,1,94.35,0,1,Offer B,3193,1,0,1,1,61,0,0.0,1533.54,29.88,5703.0,0,1,95982
6488,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.5,69.5,1,41,30,8.31,3365,1,Taylorsville,0,0,Cable,40.053684000000004,-120.74311599999999,0,72.28,0,0,None,513,0,2,0,0,1,1,0.0,8.31,0.0,69.5,0,0,95983
6489,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,18.85,18.85,1,53,0,40.49,4132,1,Twain,0,1,NA,40.022184,-121.06238400000001,0,18.85,0,0,None,73,0,1,0,0,1,5,0.0,40.49,0.0,18.85,0,0,95984
6490,1,0,0,0,26,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.4,525.55,0,29,0,6.38,4602,0,Washington,0,1,NA,39.34128,-120.78686699999999,0,19.4,0,0,None,145,0,0,0,0,26,0,0.0,165.88,4.25,525.55,1,0,95986
6491,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.2,69.2,1,44,21,23.72,4073,1,Williams,0,0,Cable,39.117537,-122.284654,0,71.968,0,0,None,4579,0,0,0,0,1,3,0.0,23.72,0.0,69.2,0,1,95987
6492,1,0,1,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.75,483.15,0,32,0,27.38,3455,0,Willows,0,1,NA,39.493990999999994,-122.286363,1,19.75,0,4,None,8812,0,0,1,0,24,0,0.0,657.12,16.56,483.15,0,0,95988
6493,1,0,1,0,17,0,No phone service,DSL,0,0,1,1,One year,0,Electronic check,54.6,934.8,0,29,27,0.0,4590,0,Yuba City,1,1,DSL,39.027409999999996,-121.61498200000001,1,54.6,0,5,Offer D,34967,1,0,1,1,17,1,252.0,0.0,47.73,934.8,1,0,95991
6494,0,0,0,1,26,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,29.8,786.5,0,24,27,0.0,3746,0,Yuba City,1,0,Cable,39.075694,-121.70606000000001,0,29.8,2,0,None,27786,0,0,0,0,26,2,21.24,0.0,10.28,786.5,1,1,95993
6495,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.65,69.65,1,30,76,28.7,5258,1,Redding,0,1,Cable,40.587919,-122.46473200000001,0,72.436,0,0,Offer E,31586,0,1,0,0,1,1,0.0,28.7,0.0,69.65,0,0,96001
6496,1,1,1,0,40,1,1,Fiber optic,1,0,1,1,Month-to-month,0,Electronic check,101.85,4086.3,1,76,3,2.85,2837,1,Redding,0,1,Fiber Optic,40.527834000000006,-122.318749,1,105.924,0,1,None,30338,0,0,1,0,40,3,12.26,114.0,0.0,4086.3,0,1,96002
6497,1,0,0,0,52,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,103.05,5364.8,0,33,22,5.42,5432,0,Redding,1,1,DSL,40.677649,-122.29467,0,103.05,0,0,Offer B,41476,0,0,0,1,52,2,1180.0,281.84,46.67,5364.8,0,0,96003
6498,0,0,0,0,1,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,82.3,82.3,1,64,31,33.41,4278,1,Adin,1,0,Cable,41.171578000000004,-120.91316100000002,0,85.59200000000001,0,0,Offer E,615,0,4,0,0,1,4,0.0,33.41,0.0,82.3,0,0,96006
6499,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.3,20.3,0,22,0,29.19,5203,0,Anderson,0,1,NA,40.448632,-122.306657,0,20.3,0,0,None,21418,0,0,0,0,1,0,0.0,29.19,0.0,20.3,1,0,96007
6500,0,0,0,0,21,0,No phone service,DSL,1,0,0,0,Two year,0,Mailed check,35.1,770.4,0,34,4,0.0,2991,0,Bella Vista,0,0,Cable,40.722733000000005,-122.10966599999999,0,35.1,0,0,Offer D,899,1,0,0,0,21,2,31.0,0.0,0.0,770.4,0,0,96008
6501,0,0,1,0,67,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),105.7,6816.95,0,23,73,25.46,5027,0,Bieber,1,0,Fiber Optic,41.083464,-121.107929,1,105.7,0,2,Offer A,595,0,0,1,1,67,1,0.0,1705.8200000000004,0.0,6816.95,1,1,96009
6502,0,0,1,1,44,1,0,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),56.25,2419.55,0,36,75,43.7,3918,0,Big Bar,0,0,DSL,40.775271999999994,-123.28741399999998,1,56.25,3,10,Offer B,269,1,0,1,0,44,0,1815.0,1922.8,14.78,2419.55,0,0,96010
6503,1,0,1,1,70,0,No phone service,DSL,0,1,1,1,One year,0,Electronic check,60.35,4138.7,0,19,47,0.0,4122,0,Big Bend,1,1,Fiber Optic,41.096569,-121.87908200000001,1,60.35,3,1,Offer A,265,1,0,1,1,70,2,1945.0,0.0,49.23,4138.7,1,0,96011
6504,1,0,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,79.25,267.6,1,33,3,49.76,4183,1,Burney,0,1,Fiber Optic,40.946785,-121.719489,0,82.42,0,0,Offer E,4552,0,1,0,0,3,4,8.0,149.28,0.0,267.6,0,0,96013
6505,1,0,1,1,56,1,0,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),59.8,3457.45,0,45,13,22.74,4964,0,Callahan,1,1,Fiber Optic,41.388397,-122.79463600000001,1,59.8,2,1,Offer B,290,0,0,1,0,56,0,0.0,1273.4399999999996,35.01,3457.45,0,1,96014
6506,0,0,0,0,13,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,84.6,1115.2,1,27,46,35.96,2659,1,Canby,0,0,Cable,41.486953,-120.913975,0,87.984,0,0,Offer D,417,0,0,0,1,13,3,513.0,467.48,0.0,1115.2,1,0,96015
6507,0,0,1,1,58,1,1,Fiber optic,1,1,0,1,Month-to-month,1,Bank transfer (automatic),93.4,5435.6,1,37,22,3.65,5989,1,Cassel,0,0,Cable,40.936285,-121.57269199999999,1,97.136,0,1,None,344,0,1,1,1,58,1,119.58,211.7,0.0,5435.6,0,1,96016
6508,0,0,1,1,42,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,94.2,4186.3,1,25,30,6.84,5458,1,Castella,0,0,Cable,41.121108,-122.33661299999999,1,97.96799999999999,0,1,None,228,0,3,1,1,42,4,1256.0,287.28,0.0,4186.3,1,0,96017
6509,1,1,1,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,25.05,25.05,1,74,20,0.0,2119,1,Shasta Lake,0,1,Cable,40.692523,-122.369876,1,26.052000000000003,0,1,Offer E,6277,0,0,1,0,1,0,0.0,0.0,0.0,25.05,0,1,96019
6510,0,0,1,1,46,1,1,Fiber optic,1,0,0,1,Two year,0,Mailed check,99.65,4630.2,0,32,18,49.26,4736,0,Chester,1,0,DSL,40.243494,-121.15473300000001,1,99.65,1,10,Offer B,2664,1,0,1,1,46,0,833.0,2265.96,9.35,4630.2,0,0,96020
6511,0,0,1,1,63,1,0,DSL,1,0,0,0,Two year,1,Bank transfer (automatic),50.65,3221.25,0,37,11,25.32,4847,0,Corning,0,0,Fiber Optic,39.913777,-122.289984,1,50.65,1,6,Offer B,13840,0,0,1,0,63,1,354.0,1595.16,37.04,3221.25,0,0,96021
6512,1,0,0,0,11,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,60.9,688.5,0,23,27,28.76,2726,0,Cottonwood,1,1,Fiber Optic,40.336392,-122.44853300000001,0,60.9,0,0,Offer D,12348,1,0,0,0,11,1,186.0,316.36,49.24,688.5,1,0,96022
6513,1,0,1,1,15,1,1,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),59.65,867.1,0,22,59,24.36,3974,0,Dorris,1,1,Fiber Optic,41.949216,-122.05006200000001,1,59.65,2,6,Offer D,1162,1,0,1,0,15,0,0.0,365.4,32.65,867.1,1,1,96023
6514,1,0,1,0,72,0,No phone service,DSL,1,1,1,1,Two year,1,Electronic check,64.7,4746.05,0,33,12,0.0,6075,0,Douglas City,1,1,Fiber Optic,40.586588,-122.903677,1,64.7,0,8,Offer A,960,1,0,1,1,72,0,0.0,0.0,0.0,4746.05,0,1,96024
6515,0,0,0,0,29,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),25.1,712.85,1,53,24,0.0,2796,1,Dunsmuir,0,0,Cable,41.212695000000004,-122.392067,0,26.104000000000006,0,0,None,2602,0,0,0,0,29,0,171.0,0.0,0.0,712.85,0,0,96025
6516,1,0,0,1,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,48.95,48.95,1,22,57,34.4,3913,1,Etna,1,1,Cable,41.405193,-123.008567,0,50.908,2,0,None,2156,0,2,0,1,1,4,0.0,34.4,0.0,48.95,1,0,96027
6517,0,0,1,1,6,1,0,DSL,0,0,1,0,Month-to-month,0,Electronic check,54.85,355.1,0,23,48,30.17,5729,0,Fall River Mills,0,0,Fiber Optic,41.017282,-121.46894499999999,1,54.85,2,3,None,1902,0,0,1,0,6,2,170.0,181.02,39.15,355.1,1,0,96028
6518,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,45.3,45.3,1,59,8,28.37,5774,1,Flournoy,0,1,Fiber Optic,39.847840000000005,-122.544556,0,47.111999999999995,0,0,None,84,0,0,0,0,1,2,0.0,28.37,0.0,45.3,0,0,96029
6519,1,0,1,1,63,1,1,Fiber optic,0,1,0,1,One year,1,Electronic check,91.35,5764.7,0,62,28,48.62,4512,0,Forks Of Salmon,0,1,Cable,41.232128,-123.194748,1,91.35,2,4,Offer B,170,0,0,1,1,63,2,1614.0,3063.06,18.78,5764.7,0,0,96031
6520,1,0,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.85,167.3,1,58,31,14.14,3273,1,Escondido,1,1,Fiber Optic,33.141265000000004,-116.967221,0,89.28399999999998,0,0,Offer E,48690,0,0,0,1,2,0,52.0,28.28,0.0,167.3,0,0,92027
6521,0,0,1,1,18,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,25.1,428.45,0,33,0,39.56,3675,0,French Gulch,0,0,NA,40.740138,-122.587476,1,25.1,1,2,Offer D,373,0,0,1,0,18,0,0.0,712.08,14.57,428.45,0,0,96033
6522,0,0,1,0,43,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),34.0,1505.35,0,34,21,0.0,5409,0,Gazelle,0,0,DSL,41.411315,-122.697236,1,34.0,0,9,Offer B,392,1,0,1,0,43,0,316.0,0.0,49.22,1505.35,0,0,96034
6523,0,0,0,0,15,0,No phone service,DSL,1,1,0,0,One year,0,Mailed check,45.9,693.45,0,60,25,0.0,3572,0,Gerber,1,0,DSL,40.031940000000006,-122.176023,0,45.9,0,0,Offer D,3357,1,0,0,0,15,2,0.0,0.0,16.27,693.45,0,1,96035
6524,1,0,0,1,10,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,95.2,930.4,1,54,20,35.63,4922,1,Greenview,0,1,DSL,41.528541,-122.955018,0,99.008,0,0,Offer D,295,0,0,0,1,10,4,18.61,356.3,0.0,930.4,0,1,96037
6525,1,0,1,1,55,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.5,1177.95,0,57,0,40.94,5011,0,Grenada,0,1,NA,41.599978,-122.539381,1,20.5,3,1,Offer B,616,0,0,1,0,55,0,0.0,2251.7,5.83,1177.95,0,0,96038
6526,1,0,0,1,49,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),100.6,5069.65,1,42,3,18.97,5585,1,Happy Camp,0,1,Cable,41.831901,-123.487478,0,104.624,0,0,None,1294,1,2,0,1,49,3,152.0,929.53,0.0,5069.65,0,0,96039
6527,1,0,1,1,6,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,55.3,324.25,1,49,21,1.86,3878,1,Hat Creek,1,1,Fiber Optic,40.789799,-121.474529,1,57.512,1,1,Offer E,397,0,1,1,0,6,2,68.0,11.16,0.0,324.25,0,0,96040
6528,1,0,1,1,70,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.35,1458.1,0,38,0,31.78,5748,0,Fallbrook,0,1,NA,33.362575,-117.299644,1,20.35,1,2,Offer A,42239,0,2,1,0,70,1,0.0,2224.6,35.44,1458.1,0,0,92028
6529,1,1,0,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.85,156.4,1,79,20,45.41,5378,1,Hornbrook,0,1,DSL,41.962127,-122.52769599999999,0,77.844,0,0,Offer E,1026,0,0,0,0,2,4,31.0,90.82,0.0,156.4,0,0,96044
6530,1,1,1,0,63,0,No phone service,DSL,1,0,0,0,One year,0,Bank transfer (automatic),36.1,2298.9,0,76,7,0.0,5089,0,Hyampom,0,1,Fiber Optic,40.648024,-123.465088,1,36.1,0,2,Offer B,268,1,0,1,0,63,0,0.0,0.0,0.0,2298.9,0,1,96046
6531,0,0,0,0,25,1,0,DSL,0,1,0,1,Month-to-month,1,Bank transfer (automatic),65.8,1679.65,0,33,10,1.22,3962,0,Igo,0,0,Fiber Optic,40.524535,-122.647172,0,65.8,0,0,None,911,1,0,0,1,25,0,168.0,30.5,29.29,1679.65,0,0,96047
6532,0,1,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.35,369.6,0,77,0,37.53,4713,0,Junction City,0,0,NA,40.913191999999995,-123.06597,0,20.35,0,0,Offer D,734,0,0,0,0,18,1,0.0,675.54,0.0,369.6,0,0,96048
6533,1,1,1,0,28,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.8,2998,0,67,15,24.35,4174,0,Klamath River,0,1,Cable,41.816595,-122.94828700000001,1,105.8,0,8,Offer C,482,1,1,1,1,28,4,450.0,681.8000000000002,0.0,2998.0,0,0,96050
6534,0,1,0,0,53,1,0,Fiber optic,1,1,0,1,One year,1,Mailed check,96.75,5206.55,0,72,28,34.58,4766,0,Lakehead,0,0,Fiber Optic,40.883853,-122.41825800000001,0,96.75,0,0,Offer B,1236,1,0,0,1,53,2,0.0,1832.74,0.0,5206.55,0,1,96051
6535,1,0,0,0,35,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),102.35,3626.1,1,26,53,39.84,2473,1,Lewiston,1,1,DSL,40.704293,-122.803899,0,106.444,0,0,None,1845,0,0,0,1,35,5,1922.0,1394.4,0.0,3626.1,1,0,96052
6536,1,0,0,0,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,24.4,24.4,0,45,29,0.0,4570,0,Lookout,0,1,DSL,41.280478,-121.160249,0,24.4,0,0,None,386,0,0,0,0,1,1,0.0,0.0,0.0,24.4,0,1,96054
6537,1,0,1,0,70,1,1,Fiber optic,1,1,1,1,One year,0,Credit card (automatic),115.65,7968.85,1,51,22,17.17,5563,1,Los Molinos,1,1,Fiber Optic,40.059385,-122.091481,1,120.276,0,1,Offer A,3756,1,0,1,1,70,0,1753.0,1201.9,0.0,7968.85,0,0,96055
6538,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,79.85,152.45,1,46,2,16.14,3280,1,Mcarthur,1,1,DSL,41.108309999999996,-121.36036200000001,0,83.044,0,0,Offer E,1554,1,1,0,0,2,3,3.0,32.28,0.0,152.45,0,0,96056
6539,0,0,1,0,26,1,0,DSL,0,1,1,1,Month-to-month,1,Electronic check,73.05,1959.5,0,35,20,23.31,2753,0,Mccloud,0,0,Fiber Optic,41.251321999999995,-122.105209,1,73.05,0,7,None,1586,1,1,1,1,26,1,0.0,606.06,47.59,1959.5,0,1,96057
6540,0,0,0,0,34,1,0,DSL,1,1,0,1,One year,0,Electronic check,64.35,2053.05,0,55,7,45.56,3445,0,Macdoel,0,0,Fiber Optic,41.769709000000006,-121.92063,0,64.35,0,0,None,816,0,0,0,1,34,0,14.37,1549.04,46.39,2053.05,0,1,96058
6541,0,0,0,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.5,398.55,0,29,0,35.45,4855,0,Manton,0,0,NA,40.426679,-121.850421,0,20.5,1,0,Offer D,598,0,0,0,0,19,1,0.0,673.5500000000002,24.07,398.55,1,0,96059
6542,1,0,0,0,15,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,76.0,1130.85,1,29,57,44.86,4938,1,Mill Creek,0,1,DSL,40.331975,-121.460674,0,79.04,0,0,Offer D,78,0,1,0,1,15,4,645.0,672.9,0.0,1130.85,1,0,96061
6543,0,0,1,1,62,1,0,DSL,1,0,0,0,One year,0,Credit card (automatic),54.75,3425.35,0,22,71,32.92,5010,0,Millville,1,0,Fiber Optic,40.531257000000004,-122.14813899999999,1,54.75,3,5,Offer B,830,0,0,1,0,62,1,0.0,2041.04,8.5,3425.35,1,1,96062
6544,0,1,0,0,42,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),104.75,4323.45,1,69,13,16.22,2984,1,Mineral,1,0,DSL,40.408796,-121.579609,0,108.94,0,0,None,124,0,2,0,0,42,1,562.0,681.24,0.0,4323.45,0,0,96063
6545,0,0,0,0,9,1,0,DSL,1,1,1,1,Month-to-month,1,Electronic check,74.65,703.55,1,31,18,36.43,5900,1,Fallbrook,0,0,DSL,33.362575,-117.299644,0,77.63600000000002,0,0,Offer E,42239,0,1,0,1,9,5,0.0,327.87,0.0,703.55,0,1,92028
6546,1,0,0,0,24,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,51.15,1275.7,0,60,22,33.97,5796,0,Montgomery Creek,0,1,DSL,40.877552,-121.885884,0,51.15,0,0,None,431,0,0,0,0,24,0,28.07,815.28,0.0,1275.7,0,1,96065
6547,1,1,1,0,68,0,No phone service,DSL,1,1,0,0,Two year,1,Electronic check,41.95,2965.75,0,79,28,0.0,5607,0,Mount Shasta,1,1,Fiber Optic,41.33832,-122.290756,1,41.95,0,9,None,7309,0,0,1,0,68,0,0.0,0.0,0.0,2965.75,0,1,96067
6548,1,0,1,1,31,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,54.35,1647,0,20,71,25.04,3615,0,Nubieber,1,1,Fiber Optic,41.082471999999996,-121.19521499999999,1,54.35,1,6,None,240,1,0,1,0,31,1,1169.0,776.24,0.0,1647.0,1,0,96068
6549,0,0,0,0,1,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,56.25,56.25,1,49,24,26.14,3065,1,Oak Run,0,0,Fiber Optic,40.689243,-122.037023,0,58.5,0,0,None,829,0,1,0,1,1,2,0.0,26.14,0.0,56.25,0,0,96069
6550,1,0,1,0,21,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,106.1,2249.95,1,27,65,21.83,3584,1,Old Station,1,1,Cable,40.656287,-121.42896499999999,1,110.344,0,1,Offer D,182,1,0,1,1,21,5,1462.0,458.43,0.0,2249.95,1,0,96071
6551,0,0,1,0,63,1,0,Fiber optic,0,1,1,1,One year,1,Electronic check,96.0,6109.75,0,20,51,20.51,5016,0,Palo Cedro,0,0,DSL,40.582399,-122.19551200000001,1,96.0,0,5,Offer B,4931,0,0,1,1,63,0,0.0,1292.13,0.0,6109.75,1,1,96073
6552,0,1,0,0,2,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),79.75,159.4,1,74,25,39.63,4038,1,Paskenta,0,0,DSL,39.884395,-122.58751299999999,0,82.94,0,0,Offer E,263,0,0,0,0,2,0,40.0,79.26,0.0,159.4,0,0,96074
6553,0,0,1,1,61,0,No phone service,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),61.45,3751.15,0,46,26,0.0,5063,0,Paynes Creek,1,0,DSL,40.343213,-121.81541200000001,1,61.45,3,8,Offer B,433,1,0,1,1,61,0,0.0,0.0,0.0,3751.15,0,1,96075
6554,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,68.65,68.65,1,62,31,12.4,3052,1,Platina,0,0,Cable,40.367964,-122.937379,0,71.39600000000002,0,0,Offer E,215,0,1,0,0,1,2,0.0,12.4,0.0,68.65,0,0,96076
6555,1,0,0,0,18,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.65,411.25,0,32,0,1.42,4695,0,Red Bluff,0,1,NA,40.186772,-122.388361,0,19.65,0,0,Offer D,26438,0,0,0,0,18,2,0.0,25.56,0.0,411.25,0,0,96080
6556,0,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.0,105.5,0,38,0,30.01,5518,0,Round Mountain,0,0,NA,40.923558,-122.059933,1,19.0,3,0,None,459,0,1,0,0,6,2,0.0,180.06,0.0,105.5,0,0,96084
6557,0,0,0,0,33,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.0,3320.6,0,44,30,16.57,4643,0,Scott Bar,0,0,Cable,41.737961999999996,-123.07557,0,100.0,0,0,None,88,0,0,0,1,33,1,996.0,546.8100000000002,0.0,3320.6,0,0,96085
6558,1,0,0,0,16,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.25,327.45,1,24,0,21.04,4327,1,Seiad Valley,0,1,NA,41.924174,-123.26078799999999,0,20.25,0,0,Offer D,332,0,2,0,0,16,4,0.0,336.64,0.0,327.45,1,0,96086
6559,0,0,1,0,56,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,98.7,5669.5,0,62,18,7.0,5141,0,Shasta,1,0,Fiber Optic,40.617614,-122.51286100000002,1,98.7,0,3,Offer B,528,1,0,1,1,56,1,0.0,392.0,0.0,5669.5,0,1,96087
6560,1,0,0,1,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.8,465.45,0,50,0,1.2,3058,0,Shingletown,0,1,NA,40.497440999999995,-121.827524,0,19.8,3,0,Offer D,4231,0,0,0,0,23,1,0.0,27.6,0.0,465.45,0,0,96088
6561,1,0,0,0,9,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,73.8,704.3,0,54,22,1.85,4895,0,Tehama,1,1,Fiber Optic,40.021786999999996,-122.127576,0,73.8,0,0,None,405,0,0,0,0,9,1,155.0,16.650000000000002,0.0,704.3,0,0,96090
6562,0,1,1,0,14,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,100.2,1369.8,1,71,21,47.01,3369,1,Trinity Center,0,0,Fiber Optic,41.081846999999996,-122.70054499999999,1,104.208,0,1,None,734,0,0,1,0,14,0,0.0,658.14,0.0,1369.8,0,1,96091
6563,1,0,1,1,15,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.9,1107.25,1,39,16,34.63,2510,1,Vina,0,1,Cable,39.955164,-122.01856699999999,1,77.89600000000002,0,1,Offer D,439,0,0,1,0,15,2,177.0,519.45,0.0,1107.25,0,0,96092
6564,1,0,0,0,5,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.05,95.55,0,26,0,22.16,2483,0,Weaverville,0,1,NA,40.759401000000004,-122.93933700000001,0,20.05,0,0,None,3749,0,1,0,0,5,2,0.0,110.8,0.0,95.55,1,0,96093
6565,1,0,1,0,61,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Electronic check,106.2,6375.2,0,40,29,27.66,6298,0,Weed,0,1,Cable,41.465121,-122.38094699999999,1,106.2,0,6,None,5896,0,0,1,1,61,0,1849.0,1687.26,0.0,6375.2,0,0,96094
6566,1,0,1,1,70,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),116.55,8152.3,0,21,71,40.77,6116,0,Whitmore,1,1,Fiber Optic,40.637105,-121.906949,1,116.55,2,5,Offer A,843,1,0,1,1,70,1,5788.0,2853.9,0.0,8152.3,1,0,96096
6567,1,0,0,0,15,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,99.7,1566.75,0,53,15,10.12,4157,0,Yreka,0,1,DSL,41.764869,-122.67131599999999,0,99.7,0,0,Offer D,9538,0,0,0,1,15,0,23.5,151.79999999999995,0.0,1566.75,0,1,96097
6568,1,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.7,130.25,0,27,0,11.57,5962,0,Alturas,0,1,NA,41.468877,-120.54229,1,19.7,1,8,None,5096,0,0,1,0,8,2,0.0,92.56,0.0,130.25,1,0,96101
6569,0,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.5,162.15,0,19,0,13.21,3598,0,Blairsden Graeagle,0,0,NA,39.783747,-120.661032,1,19.5,2,10,None,1839,0,0,1,0,8,0,0.0,105.68,0.0,162.15,1,0,96103
6570,0,0,0,0,4,0,No phone service,DSL,1,0,0,0,Month-to-month,1,Mailed check,29.15,110.05,0,53,2,0.0,2657,0,Cedarville,0,0,Cable,41.505916,-120.152505,0,29.15,0,0,None,857,0,0,0,0,4,1,0.0,0.0,0.0,110.05,0,1,96104
6571,0,0,0,0,34,1,0,DSL,1,1,0,0,One year,0,Mailed check,55.0,1885.15,0,31,8,43.17,4027,0,Chilcoot,0,0,DSL,39.872961,-120.198876,0,55.0,0,0,Offer C,650,0,0,0,0,34,0,151.0,1467.78,0.0,1885.15,0,0,96105
6572,1,0,1,0,68,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),90.8,6302.85,0,38,21,11.83,4265,0,Clio,1,1,Fiber Optic,39.745805,-120.580882,1,90.8,0,1,Offer A,88,1,0,1,1,68,0,0.0,804.44,0.0,6302.85,0,1,96106
6573,0,0,1,1,45,0,No phone service,DSL,0,1,0,1,One year,0,Bank transfer (automatic),51.0,2264.5,0,52,19,0.0,4534,0,Coleville,1,0,Cable,38.42528,-119.47574099999999,1,51.0,2,10,None,1332,1,0,1,1,45,2,43.03,0.0,0.0,2264.5,0,1,96107
6574,0,1,0,0,9,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,90.1,816.8,0,66,4,40.0,2893,0,Davis Creek,1,0,Fiber Optic,41.750353999999994,-120.403885,0,90.1,0,0,Offer E,104,0,0,0,0,9,0,0.0,360.0,0.0,816.8,0,1,96108
6575,0,0,0,0,22,1,1,DSL,1,0,0,0,Month-to-month,1,Mailed check,59.05,1253.5,0,33,24,32.75,3995,0,Doyle,0,0,DSL,40.012675,-120.10185700000001,0,59.05,0,0,Offer D,1177,1,0,0,0,22,0,0.0,720.5,0.0,1253.5,0,1,96109
6576,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.3,41.2,0,39,0,12.68,5074,0,Eagleville,0,0,NA,41.280341,-120.15038100000001,0,20.3,0,0,None,132,0,2,0,0,2,2,0.0,25.36,0.0,41.2,0,0,96110
6577,1,0,1,0,70,1,1,DSL,0,1,1,0,Two year,0,Bank transfer (automatic),72.95,5265.55,0,50,25,38.58,6466,0,Fort Bidwell,1,1,Cable,41.932207,-120.13594099999999,1,72.95,0,4,Offer A,231,1,0,1,0,70,0,0.0,2700.6,0.0,5265.55,0,1,96112
6578,0,0,0,1,10,1,1,DSL,1,0,0,1,One year,0,Credit card (automatic),73.55,693.3,0,23,26,14.24,4434,0,Herlong,1,0,Fiber Optic,40.198234,-120.18088999999999,0,73.55,1,0,Offer D,946,1,1,0,1,10,2,0.0,142.4,0.0,693.3,1,1,96113
6579,1,0,0,0,72,1,1,DSL,1,0,1,1,Two year,0,Credit card (automatic),84.3,5997.1,0,55,27,29.03,6012,0,Janesville,1,1,DSL,40.294034,-120.512622,0,84.3,0,0,Offer A,3093,1,1,0,1,72,1,1619.0,2090.16,0.0,5997.1,0,0,96114
6580,0,0,1,1,49,1,0,DSL,0,1,1,1,One year,0,Credit card (automatic),78.0,3824.2,0,23,82,9.07,4200,0,Fallbrook,1,0,Fiber Optic,33.362575,-117.299644,1,78.0,1,10,None,42239,0,0,1,1,49,0,0.0,444.43,0.0,3824.2,1,1,92028
6581,0,1,0,0,54,1,1,DSL,0,1,1,0,One year,0,Mailed check,72.1,3886.05,0,68,2,45.43,4277,0,Likely,0,0,Fiber Optic,41.266008,-120.49073100000001,0,72.1,0,0,Offer B,277,1,0,0,0,54,0,7.77,2453.22,0.0,3886.05,0,1,96116
6582,0,0,0,0,71,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),106.75,7283.25,0,57,10,2.93,5610,0,Litchfield,1,0,Fiber Optic,40.507272,-120.338228,0,106.75,0,0,Offer A,385,0,0,0,1,71,0,0.0,208.03,0.0,7283.25,0,1,96117
6583,0,0,0,0,22,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.25,412.55,0,50,0,35.4,2691,0,Loyalton,0,0,NA,39.637471000000005,-120.22633799999998,0,19.25,0,0,None,1822,0,0,0,0,22,1,0.0,778.8,0.0,412.55,0,0,96118
6584,0,0,1,1,50,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.55,1070.25,0,37,0,10.13,4878,0,Madeline,0,0,NA,41.042003,-120.50608600000001,1,20.55,3,10,None,85,0,0,1,0,50,2,0.0,506.50000000000006,0.0,1070.25,0,0,96119
6585,0,0,1,1,43,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.0,817.95,0,51,0,35.2,4882,0,Markleeville,0,0,NA,38.735789000000004,-119.85798,1,20.0,2,5,None,957,0,0,1,0,43,2,0.0,1513.6,0.0,817.95,0,0,96120
6586,0,0,1,1,45,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),24.65,1171.3,0,21,0,37.57,2194,0,Milford,0,0,NA,40.181278999999996,-120.392967,1,24.65,1,5,None,481,0,0,1,0,45,1,0.0,1690.65,0.0,1171.3,1,0,96121
6587,1,1,0,0,64,1,1,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),103.5,6548.65,0,78,18,19.2,5125,0,Portola,0,1,Fiber Optic,39.786755,-120.445626,0,103.5,0,0,Offer B,4236,0,0,0,1,64,0,0.0,1228.8,0.0,6548.65,0,1,96122
6588,0,0,1,1,23,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,23.85,625.65,0,61,0,7.11,5945,0,Ravendale,0,0,NA,40.845738,-120.32221899999999,1,23.85,3,0,None,61,0,0,0,0,23,0,0.0,163.53,0.0,625.65,0,0,96123
6589,0,0,1,0,68,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.8,1911.5,0,41,0,17.12,4747,0,Calpine,0,0,NA,39.672813,-120.456699,1,25.8,0,8,Offer A,322,0,2,1,0,68,2,0.0,1164.16,0.0,1911.5,0,0,96124
6590,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.85,70.85,1,51,25,27.05,2874,1,Sierra City,0,0,Fiber Optic,39.600599,-120.636358,0,73.684,0,0,Offer E,348,0,3,0,0,1,3,0.0,27.05,0.0,70.85,0,1,96125
6591,1,0,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),69.8,134.7,1,56,30,37.72,2320,1,Sierraville,0,1,Cable,39.559709000000005,-120.34563899999999,0,72.592,0,0,Offer E,227,0,1,0,0,2,3,40.0,75.44,0.0,134.7,0,0,96126
6592,1,0,0,0,26,1,0,DSL,0,0,1,0,One year,0,Credit card (automatic),59.45,1507,0,47,6,3.26,2074,0,Standish,0,1,DSL,40.346634,-120.386422,0,59.45,0,0,Offer C,408,1,0,0,0,26,0,0.0,84.75999999999998,0.0,1507.0,0,1,96128
6593,1,0,1,0,55,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Bank transfer (automatic),54.55,2978.3,1,30,46,0.0,6041,1,Susanville,1,1,Fiber Optic,40.559177000000005,-120.612113,1,56.732,0,1,None,19440,1,0,1,1,55,2,1370.0,0.0,0.0,2978.3,0,0,96130
6594,1,0,0,0,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.05,299.3,0,27,0,9.19,5728,0,Termo,0,1,NA,41.027281,-120.669427,0,20.05,0,0,None,72,0,0,0,0,14,0,0.0,128.66,0.0,299.3,1,0,96132
6595,1,0,1,0,71,1,0,DSL,1,0,1,1,Two year,1,Electronic check,82.55,5832.65,0,34,19,28.21,4668,0,Topaz,1,1,DSL,38.636052,-119.48916200000001,1,82.55,0,2,Offer A,116,1,0,1,1,71,3,0.0,2002.91,0.0,5832.65,0,1,96133
6596,1,0,0,0,64,1,1,DSL,1,1,1,0,One year,0,Electronic check,81.25,5567.55,0,25,69,5.49,4761,0,Tulelake,1,1,DSL,41.813521,-121.49266599999999,0,81.25,0,0,None,2595,1,0,0,0,64,0,0.0,351.36,0.0,5567.55,1,1,96134
6597,0,0,0,0,7,1,0,DSL,0,0,1,1,Month-to-month,1,Credit card (automatic),70.75,450.8,1,57,7,23.35,2248,1,Wendel,0,0,Cable,40.345949,-120.08118700000001,0,73.58,0,0,Offer E,162,1,2,0,1,7,3,32.0,163.45000000000005,0.0,450.8,0,0,96136
6598,0,0,0,0,57,1,0,DSL,1,1,1,0,Two year,1,Credit card (automatic),74.3,4166.35,0,61,3,6.45,5741,0,Westwood,1,0,Fiber Optic,40.271535,-121.01808700000001,0,74.3,0,0,None,4158,1,0,0,0,57,2,0.0,367.65,0.0,4166.35,0,1,96137
6599,0,0,1,0,13,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Electronic check,94.1,1215.6,1,26,57,43.56,2973,1,Carnelian Bay,1,0,Cable,39.227434,-120.091806,1,97.86399999999999,0,1,None,1943,0,1,1,0,13,3,693.0,566.28,0.0,1215.6,1,0,96140
6600,0,0,1,1,3,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),29.7,91.7,1,46,16,0.0,2613,1,Homewood,0,0,DSL,39.117018,-120.212535,1,30.888,2,1,Offer E,858,0,0,1,0,3,5,15.0,0.0,0.0,91.7,0,0,96141
6601,1,1,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,0,Credit card (automatic),109.7,7898.45,0,76,3,27.74,4319,0,Tahoma,1,1,Fiber Optic,39.061227,-120.179546,1,109.7,0,5,None,1291,1,0,1,1,72,0,0.0,1997.28,0.0,7898.45,0,1,96142
6602,0,0,1,1,40,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),96.35,3915.4,0,51,23,29.42,2004,0,Kings Beach,1,0,Fiber Optic,39.246654,-120.029273,1,96.35,2,4,None,4806,0,0,1,0,40,1,0.0,1176.8000000000004,0.0,3915.4,0,1,96143
6603,1,0,1,0,14,1,1,DSL,0,0,1,0,Month-to-month,1,Credit card (automatic),66.6,979.5,0,48,11,22.14,3516,0,Tahoe City,0,1,DSL,39.178337,-120.162806,1,66.6,0,3,None,4002,1,0,1,0,14,2,108.0,309.9600000000001,0.0,979.5,0,0,96145
6604,1,0,1,1,2,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,44.5,90.05,0,33,19,30.87,5456,0,Olympic Valley,0,1,Fiber Optic,39.191796999999994,-120.212401,1,44.5,1,2,None,942,0,0,1,0,2,1,0.0,61.74,0.0,90.05,0,1,96146
6605,1,1,0,0,66,1,1,Fiber optic,0,1,1,1,One year,0,Credit card (automatic),110.9,7432.05,1,69,28,9.9,4389,1,Tahoe Vista,1,1,Cable,39.241240000000005,-120.05476499999999,0,115.336,0,0,None,678,1,0,0,0,66,2,2081.0,653.4,0.0,7432.05,0,0,96148
6606,0,0,1,0,38,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,105.0,4026.4,1,60,4,19.08,2341,1,San Diego,1,0,Fiber Optic,32.898613,-117.202937,1,109.2,0,1,None,4258,1,0,1,1,38,1,161.0,725.04,0.0,4026.4,0,0,92121
6607,1,0,0,1,1,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,25.3,25.3,1,20,56,0.0,5421,1,San Diego,0,1,Cable,32.898613,-117.202937,0,26.311999999999998,3,0,None,4258,0,2,0,0,1,3,0.0,0.0,0.0,25.3,1,0,92121
6608,1,0,0,0,22,1,0,DSL,0,1,0,0,One year,1,Credit card (automatic),55.15,1193.05,1,22,65,33.53,5866,1,San Diego,0,1,Cable,32.898613,-117.202937,0,57.356,0,0,None,4258,1,2,0,0,22,5,775.0,737.6600000000002,0.0,1193.05,1,0,92121
6609,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.1,20.1,1,25,0,4.11,4389,1,San Diego,0,1,NA,32.898613,-117.202937,0,20.1,0,0,None,4258,0,1,0,0,1,4,0.0,4.11,0.0,20.1,1,0,92121
6610,1,0,0,0,5,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,80.1,398.55,0,56,13,12.35,5225,0,Los Angeles,0,1,Cable,33.964131,-118.272783,0,80.1,0,0,None,58198,0,0,0,0,5,2,0.0,61.75,0.0,398.55,0,1,90003
6611,1,0,1,1,29,1,1,DSL,1,0,1,0,One year,0,Bank transfer (automatic),69.05,1958.45,0,26,69,36.7,4459,0,Los Angeles,0,1,DSL,34.076259,-118.31071499999999,1,69.05,2,5,Offer C,67852,1,0,1,0,29,2,135.13,1064.3000000000004,0.0,1958.45,1,1,90004
6612,1,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.9,69.9,1,49,31,4.99,2100,1,San Diego,0,1,Cable,32.898613,-117.202937,1,72.69600000000001,0,0,None,4258,0,0,0,0,1,4,0.0,4.99,0.0,69.9,0,0,92121
6613,0,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.4,63.15,0,42,0,14.79,5695,0,Los Angeles,0,0,NA,34.048013,-118.293953,0,20.4,0,0,Offer E,62784,0,0,0,0,3,1,0.0,44.37,0.0,63.15,0,0,90006
6614,1,0,1,1,71,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.7,1301.1,0,53,0,14.86,4808,0,Los Angeles,0,1,NA,34.027337,-118.28515,1,19.7,1,8,Offer A,45025,0,0,1,0,71,2,0.0,1055.06,0.0,1301.1,0,0,90007
6615,1,0,0,1,9,1,0,DSL,0,1,0,0,Month-to-month,1,Electronic check,50.1,484.05,0,34,29,27.64,4738,0,Los Angeles,0,1,Cable,34.008293,-118.34676599999999,0,50.1,2,0,Offer E,30852,0,0,0,0,9,1,14.04,248.76,0.0,484.05,0,1,90008
6616,1,0,0,0,43,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,101.4,4528,1,39,30,49.64,3370,1,San Diego,0,1,Fiber Optic,32.898613,-117.202937,0,105.456,0,0,None,4258,0,1,0,1,43,2,1358.0,2134.52,0.0,4528.0,0,0,92121
6617,0,0,0,0,48,1,1,DSL,1,1,1,1,One year,1,Credit card (automatic),83.45,3887.85,0,30,27,45.51,4250,0,Los Angeles,1,0,Fiber Optic,34.007090000000005,-118.25868100000001,0,83.45,0,0,None,101215,0,0,0,1,48,0,104.97,2184.48,0.0,3887.85,0,1,90011
6618,1,0,0,0,26,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),86.65,2208.75,0,19,48,49.87,4469,0,Los Angeles,0,1,DSL,34.065875,-118.23872800000001,0,86.65,0,0,Offer C,30596,0,0,0,0,26,0,106.02,1296.62,0.0,2208.75,1,1,90012
6619,0,0,0,0,9,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),20.15,238.15,0,63,0,34.79,3772,0,Los Angeles,0,0,NA,34.044639000000004,-118.24041299999999,0,20.15,0,0,Offer E,9732,0,2,0,0,9,1,0.0,313.11,0.0,238.15,0,0,90013
6620,1,0,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.8,80.8,1,34,16,41.77,4424,1,San Diego,0,1,Fiber Optic,32.898613,-117.202937,0,84.03200000000001,0,0,None,4258,0,0,0,1,1,3,0.0,41.77,0.0,80.8,0,1,92121
6621,0,0,1,1,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.4,958.15,0,46,0,12.68,4630,0,Los Angeles,0,0,NA,34.039224,-118.26629299999999,1,19.4,3,9,None,15140,0,0,1,0,46,0,0.0,583.28,0.0,958.15,0,0,90015
6622,1,0,0,0,2,1,1,DSL,0,0,0,1,Month-to-month,0,Bank transfer (automatic),62.05,118.3,1,44,22,37.29,5344,1,San Diego,0,1,DSL,32.898613,-117.202937,0,64.532,0,0,None,4258,0,0,0,1,2,1,26.0,74.58,0.0,118.3,0,0,92121
6623,1,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,76.45,76.45,1,74,14,3.84,3763,1,San Diego,0,1,DSL,32.898613,-117.202937,0,79.50800000000002,0,0,None,4258,0,0,0,0,1,6,0.0,3.84,0.0,76.45,0,0,92121
6624,1,0,1,1,64,0,No phone service,DSL,1,0,1,1,Two year,1,Bank transfer (automatic),60.05,3845.45,0,48,19,0.0,4120,0,Los Angeles,1,1,Fiber Optic,34.028735,-118.31723600000001,1,60.05,1,3,None,47143,1,0,1,1,64,0,0.0,0.0,0.0,3845.45,0,1,90018
6625,0,1,0,0,12,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,91.3,1094.5,1,79,20,34.01,4703,1,San Diego,0,0,Cable,32.898613,-117.202937,0,94.95200000000001,0,0,None,4258,0,0,0,0,12,5,219.0,408.12,0.0,1094.5,0,0,92121
6626,1,1,1,0,6,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.75,573.75,1,69,7,47.9,5750,1,San Diego,1,1,Cable,32.898613,-117.202937,1,99.58,0,0,Offer E,4258,0,0,0,0,6,3,0.0,287.4,0.0,573.75,0,1,92121
6627,0,0,1,0,59,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.35,1267,0,29,0,31.43,5757,0,Los Angeles,0,0,NA,34.029043,-118.23950400000001,1,20.35,0,6,None,3012,0,0,1,0,59,2,0.0,1854.37,0.0,1267.0,1,0,90021
6628,0,0,0,0,7,1,0,Fiber optic,0,1,1,1,One year,1,Mailed check,94.05,633.45,0,20,42,36.49,5545,0,Los Angeles,0,0,Fiber Optic,34.02381,-118.156582,0,94.05,0,0,Offer E,68701,0,0,0,1,7,0,266.0,255.43,0.0,633.45,1,0,90022
6629,0,1,1,0,72,1,1,DSL,1,1,1,1,Two year,1,Credit card (automatic),84.1,6129.65,0,72,28,47.4,4999,0,Los Angeles,1,0,DSL,34.017697,-118.200577,1,84.1,0,5,None,47487,0,0,1,1,72,0,0.0,3412.8,0.0,6129.65,0,1,90023
6630,1,1,0,0,16,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,78.75,1218.25,0,68,17,39.52,4351,0,Los Angeles,0,1,DSL,34.066303000000005,-118.435479,0,78.75,0,0,Offer D,44150,0,0,0,1,16,1,0.0,632.32,0.0,1218.25,0,1,90024
6631,1,0,1,0,25,1,1,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),55.55,1405.3,0,49,10,11.6,2950,0,Los Angeles,1,1,Fiber Optic,34.046174,-118.44633300000001,1,55.55,0,7,Offer C,41175,0,0,1,0,25,2,0.0,290.0,0.0,1405.3,0,1,90025
6632,0,0,1,0,34,1,1,DSL,1,1,0,0,Month-to-month,0,Electronic check,62.65,2274.9,1,19,78,41.32,3918,1,Los Angeles,0,0,DSL,34.078990999999995,-118.26380400000001,1,65.156,0,1,None,73686,1,1,1,0,34,3,1774.0,1404.88,0.0,2274.9,1,0,90026
6633,0,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.5,74.5,1,33,28,13.61,2016,1,Los Angeles,0,0,Fiber Optic,34.127194,-118.295647,0,77.48,0,0,None,48727,0,2,0,0,1,1,0.0,13.61,0.0,74.5,0,0,90027
6634,0,0,1,1,10,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),102.1,1068.85,1,31,24,32.07,3596,1,Los Angeles,1,0,Cable,34.099869,-118.326843,1,106.184,0,1,None,30568,0,1,1,1,10,3,257.0,320.7,0.0,1068.85,0,0,90028
6635,1,0,1,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,20.1,533.9,0,56,0,35.8,5689,0,Los Angeles,0,1,NA,34.089953,-118.294824,1,20.1,0,9,Offer C,41713,0,0,1,0,24,2,0.0,859.1999999999998,0.0,533.9,0,0,90029
6636,0,0,1,1,10,1,1,DSL,1,1,1,0,One year,0,Electronic check,70.3,676.15,0,42,26,26.37,5496,0,Los Angeles,0,0,Fiber Optic,34.085807,-118.206617,1,70.3,1,5,None,38415,0,0,1,0,10,0,17.58,263.7,0.0,676.15,0,1,90031
6637,1,0,1,0,69,1,0,DSL,1,1,0,0,One year,1,Credit card (automatic),53.65,3804.4,0,36,16,14.18,6092,0,Los Angeles,0,1,Fiber Optic,34.078821000000005,-118.177576,1,53.65,0,7,Offer A,46960,0,0,1,0,69,1,609.0,978.42,0.0,3804.4,0,0,90032
6638,1,0,0,0,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.75,1118.8,0,37,0,38.73,6271,0,Los Angeles,0,1,NA,34.050197999999995,-118.21094599999999,0,20.75,0,0,None,49431,0,0,0,0,57,1,0.0,2207.61,0.0,1118.8,0,0,90033
6639,1,0,1,1,50,1,0,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),103.4,5236.4,0,38,22,36.21,5437,0,Los Angeles,1,1,Cable,34.030578000000006,-118.39961299999999,1,103.4,1,2,None,58218,1,0,1,1,50,2,0.0,1810.5,0.0,5236.4,0,1,90034
6640,1,0,1,1,28,0,No phone service,DSL,1,0,1,0,One year,0,Mailed check,50.8,1386.8,0,42,19,0.0,3240,0,Los Angeles,1,1,DSL,34.051809000000006,-118.383843,1,50.8,1,2,Offer C,27799,1,0,1,0,28,2,0.0,0.0,0.0,1386.8,0,1,90035
6641,0,0,0,0,16,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,50.15,762.25,1,21,58,14.26,4254,1,Los Angeles,0,0,Cable,34.070291,-118.34919099999999,0,52.156000000000006,0,0,None,32901,0,0,0,0,16,2,442.0,228.16,0.0,762.25,1,0,90036
6642,1,0,0,0,25,1,0,DSL,1,1,1,1,Month-to-month,1,Mailed check,79.0,1902,0,28,71,7.55,5263,0,Los Angeles,0,1,Fiber Optic,34.002642,-118.287596,0,79.0,0,0,Offer C,56709,1,0,0,1,25,1,1350.0,188.75,0.0,1902.0,1,0,90037
6643,0,1,1,0,3,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),74.6,239.05,0,80,17,39.51,3711,0,Los Angeles,0,0,Fiber Optic,34.088017,-118.327168,1,74.6,0,3,Offer E,32562,0,0,1,0,3,0,41.0,118.53,0.0,239.05,0,0,90038
6644,1,0,1,0,61,1,1,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),96.5,5673.7,0,46,2,21.96,5926,0,Los Angeles,0,1,Fiber Optic,34.110845,-118.25959499999999,1,96.5,0,1,None,29310,0,0,1,1,61,2,113.0,1339.56,0.0,5673.7,0,0,90039
6645,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.1,39.8,0,60,0,35.5,2051,0,Los Angeles,0,0,NA,33.994524,-118.149953,0,20.1,0,0,None,9805,0,0,0,0,2,1,0.0,71.0,0.0,39.8,0,0,90040
6646,1,0,1,1,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.4,997.75,0,38,0,37.63,4025,0,Los Angeles,0,1,NA,34.137412,-118.20760700000001,1,19.4,3,3,None,27866,0,0,1,0,51,1,0.0,1919.13,0.0,997.75,0,0,90041
6647,0,0,1,1,71,1,0,DSL,1,0,1,1,Two year,0,Credit card (automatic),77.55,5574.35,0,21,71,48.76,5097,0,Los Angeles,1,0,Cable,34.11572,-118.19275400000001,1,77.55,3,10,Offer A,64672,0,0,1,1,71,0,0.0,3461.96,0.0,5574.35,1,1,90042
6648,0,0,1,1,20,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.05,406.05,0,31,0,14.79,2698,0,Los Angeles,0,0,NA,33.988543,-118.33408100000001,1,20.05,2,10,None,44764,0,0,1,0,20,0,0.0,295.7999999999999,0.0,406.05,0,0,90043
6649,1,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),19.85,138.85,0,54,0,23.73,2186,0,Los Angeles,0,1,NA,33.952714,-118.292061,1,19.85,2,8,Offer E,87383,0,0,1,0,6,0,0.0,142.38,0.0,138.85,0,0,90044
6650,0,0,0,0,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.2,123.65,0,64,0,43.18,5029,0,Los Angeles,0,0,NA,33.954017,-118.402447,0,20.2,0,0,Offer E,39334,0,0,0,0,6,1,0.0,259.08,0.0,123.65,0,0,90045
6651,0,0,0,0,29,1,1,DSL,1,1,0,0,Month-to-month,0,Mailed check,67.45,1801.1,0,48,2,13.74,3152,0,Los Angeles,0,0,DSL,34.108455,-118.362081,0,67.45,0,0,Offer C,49839,1,0,0,0,29,0,0.0,398.46,0.0,1801.1,0,1,90046
6652,1,0,0,0,36,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),18.55,689,0,33,0,8.5,5703,0,Los Angeles,0,1,NA,33.958149,-118.30844099999999,0,18.55,0,0,Offer C,47107,0,0,0,0,36,2,0.0,306.0,0.0,689.0,0,0,90047
6653,0,0,0,0,28,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,29.75,790.7,0,35,14,0.0,5463,0,Los Angeles,1,0,Cable,34.072945000000004,-118.37267,0,29.75,0,0,Offer C,21739,0,0,0,0,28,1,111.0,0.0,0.0,790.7,0,0,90048
6654,0,0,1,0,7,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.5,582.5,1,62,12,22.61,3887,1,Los Angeles,0,0,Cable,34.091829,-118.491244,1,89.96000000000002,0,1,None,33523,0,3,1,0,7,4,70.0,158.26999999999995,0.0,582.5,0,0,90049
6655,0,0,0,0,63,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,24.2,1618.2,0,64,0,26.74,4948,0,Los Angeles,0,0,NA,33.987945,-118.370442,0,24.2,0,0,Offer B,8115,0,1,0,0,63,3,0.0,1684.62,0.0,1618.2,0,0,90056
6656,1,0,1,1,48,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,23.55,1173.35,0,39,0,11.86,5019,0,Los Angeles,0,1,NA,34.061918,-118.27793899999999,1,23.55,1,0,Offer B,44004,0,0,0,0,48,1,0.0,569.28,0.0,1173.35,0,0,90057
6657,0,0,1,0,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Bank transfer (automatic),20.45,900.9,0,48,0,49.58,6061,0,Los Angeles,0,0,NA,34.001616999999996,-118.222274,1,20.45,0,5,Offer B,3642,0,0,1,0,49,0,0.0,2429.42,0.0,900.9,0,0,90058
6658,1,1,0,0,27,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,81.45,2122.05,1,80,6,42.91,2571,1,Los Angeles,0,1,Fiber Optic,33.927254,-118.249826,0,84.70800000000001,0,0,None,38128,0,0,0,0,27,6,127.0,1158.57,0.0,2122.05,0,0,90059
6659,1,0,1,0,72,1,1,DSL,1,1,1,1,Two year,0,Credit card (automatic),92.3,6719.9,0,42,5,13.59,5136,0,Los Angeles,1,1,Cable,33.921279999999996,-118.27418600000001,1,92.3,0,5,Offer A,24511,1,0,1,1,72,2,336.0,978.48,0.0,6719.9,0,0,90061
6660,1,0,1,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.15,69.15,1,54,33,2.2,4179,1,Los Angeles,0,1,DSL,34.003553000000004,-118.30893300000001,1,71.91600000000003,0,1,None,29299,0,0,1,0,1,2,0.0,2.2,0.0,69.15,0,0,90062
6661,0,0,1,1,72,0,No phone service,DSL,0,1,1,1,Two year,0,Credit card (automatic),53.65,3784,0,49,53,0.0,5498,0,Los Angeles,0,0,Cable,34.044271,-118.18523700000001,1,53.65,3,9,None,55668,1,0,1,1,72,2,0.0,0.0,0.0,3784.0,0,1,90063
6662,0,0,0,0,47,0,No phone service,DSL,1,1,0,0,One year,0,Credit card (automatic),39.65,1798.65,0,57,3,0.0,4670,0,Los Angeles,0,0,Cable,34.037251,-118.423573,0,39.65,0,0,Offer B,24505,1,0,0,0,47,1,0.0,0.0,0.0,1798.65,0,1,90064
6663,0,0,0,0,1,1,0,DSL,0,0,1,0,Month-to-month,1,Electronic check,54.65,54.65,0,41,4,36.33,5882,0,Los Angeles,0,0,Fiber Optic,34.108833000000004,-118.22971499999998,0,54.65,0,0,None,47534,0,0,0,0,1,0,0.0,36.33,0.0,54.65,0,0,90065
6664,0,0,0,0,36,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),104.8,3886.45,0,52,4,28.41,5319,0,Los Angeles,1,0,DSL,34.002028,-118.430656,0,104.8,0,0,Offer C,55204,0,0,0,1,36,2,15.55,1022.76,0.0,3886.45,0,1,90066
6665,1,0,1,1,43,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Credit card (automatic),29.3,1224.05,0,44,53,0.0,4741,0,Los Angeles,0,1,Fiber Optic,34.057496,-118.413959,1,29.3,3,5,Offer B,2527,0,0,1,0,43,0,0.0,0.0,0.0,1224.05,0,1,90067
6666,0,1,1,0,27,1,1,DSL,0,1,1,1,Month-to-month,0,Electronic check,83.85,2310.2,0,76,21,3.43,5907,0,Los Angeles,1,0,DSL,34.137411,-118.328915,1,83.85,0,5,Offer C,21728,1,0,1,1,27,0,0.0,92.61,0.0,2310.2,0,1,90068
6667,0,0,0,0,9,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,79.55,723.4,1,40,25,45.41,3246,1,West Hollywood,0,0,DSL,34.093781,-118.38106100000002,0,82.73200000000001,0,0,None,20408,0,0,0,1,9,2,181.0,408.69,0.0,723.4,0,0,90069
6668,0,0,0,0,38,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,103.65,3988.5,0,22,27,23.95,2511,0,Los Angeles,1,0,Fiber Optic,34.052917,-118.255178,0,103.65,0,0,Offer C,21,1,0,0,1,38,0,0.0,910.1,0.0,3988.5,1,1,90071
6669,0,1,0,0,35,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,99.05,3554.6,0,78,7,31.64,3484,0,Los Angeles,0,0,Cable,34.102084000000005,-118.451629,0,99.05,0,0,Offer C,10470,0,0,0,1,35,1,24.88,1107.4,0.0,3554.6,0,1,90077
6670,0,0,1,1,0,1,1,DSL,0,1,1,0,Two year,0,Mailed check,73.35, ,0,25,59,5.59,2342,0,Bell,1,0,Fiber Optic,33.970343,-118.17136799999999,1,73.35,3,6,Offer E,105285,1,0,1,0,10,2,433.0,55.9,0.0,733.5,1,0,90201
6671,0,0,1,0,59,1,0,Fiber optic,0,1,1,1,Two year,1,Mailed check,100.05,6034.85,0,32,11,45.75,4521,0,Beverly Hills,0,0,Fiber Optic,34.099891,-118.41433799999999,1,100.05,0,10,Offer B,21397,1,0,1,1,59,1,0.0,2699.25,0.0,6034.85,0,1,90210
6672,1,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.35,531.6,0,42,0,39.77,4962,0,Beverly Hills,0,1,NA,34.063947,-118.38300100000001,0,20.35,0,0,Offer C,8321,0,0,0,0,27,0,0.0,1073.7900000000004,0.0,531.6,0,0,90211
6673,0,1,0,0,2,1,0,DSL,0,0,0,0,Month-to-month,0,Electronic check,43.95,85.1,0,74,30,19.09,4057,0,Beverly Hills,0,0,DSL,34.062095,-118.401508,0,43.95,0,0,Offer E,11355,0,0,0,0,2,2,0.0,38.18,0.0,85.1,0,1,90212
6674,1,0,0,0,7,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,23.5,173,0,54,0,1.41,5508,0,Compton,0,1,NA,33.88151,-118.234451,0,23.5,0,0,Offer E,47305,0,0,0,0,7,1,0.0,9.87,0.0,173.0,0,0,90220
6675,0,0,0,0,36,1,1,DSL,0,1,0,1,One year,1,Mailed check,70.7,2511.95,0,55,9,29.27,3566,0,Compton,0,0,DSL,33.885811,-118.20645900000001,0,70.7,0,0,Offer C,51387,1,1,0,1,36,2,0.0,1053.72,0.0,2511.95,0,1,90221
6676,0,0,1,1,41,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Bank transfer (automatic),94.3,3893.6,0,19,59,1.6,2196,0,Compton,0,0,Cable,33.912246,-118.236773,1,94.3,2,10,Offer B,29825,0,0,1,0,41,0,0.0,65.60000000000001,0.0,3893.6,1,1,90222
6677,0,0,0,0,13,0,No phone service,DSL,0,1,0,0,Month-to-month,0,Electronic check,29.15,357.15,0,33,28,0.0,2876,0,Culver City,0,0,Fiber Optic,33.993990999999994,-118.39703999999999,0,29.15,0,0,None,31963,0,0,0,0,13,1,100.0,0.0,0.0,357.15,0,0,90230
6678,1,0,0,1,19,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),20.85,467.5,0,62,0,36.16,2654,0,Culver City,0,1,NA,34.019323,-118.391902,0,20.85,2,0,None,15195,0,0,0,0,19,1,0.0,687.04,0.0,467.5,0,0,90232
6679,0,0,1,0,60,0,No phone service,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),37.7,2288.7,0,61,2,0.0,5148,0,Downey,0,0,Fiber Optic,33.956228,-118.120993,1,37.7,0,1,Offer B,24908,1,0,1,0,60,2,0.0,0.0,0.0,2288.7,0,1,90240
6680,0,0,0,1,48,1,0,Fiber optic,0,1,1,0,Two year,1,Mailed check,95.5,4627.85,1,47,32,29.54,2459,1,Downey,1,0,Cable,33.940884000000004,-118.128628,0,99.32,0,0,None,40152,1,0,0,0,48,1,0.0,1417.92,0.0,4627.85,0,1,90241
6681,1,1,0,0,3,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,91.05,289.1,1,65,9,26.32,2194,1,Downey,1,1,Cable,33.921793,-118.140588,0,94.692,0,0,Offer E,42459,0,0,0,0,3,3,26.0,78.96000000000002,0.0,289.1,0,0,90242
6682,1,0,1,0,69,1,1,Fiber optic,0,1,1,0,Two year,1,Mailed check,92.45,6460.55,0,47,20,3.08,4452,0,El Segundo,0,1,Fiber Optic,33.917145,-118.401554,1,92.45,0,9,None,16041,1,0,1,0,69,2,0.0,212.52,0.0,6460.55,0,1,90245
6683,1,0,0,0,43,0,No phone service,DSL,0,0,0,1,One year,0,Electronic check,44.15,1931.3,0,63,11,0.0,2522,0,Gardena,1,1,DSL,33.890853,-118.29796699999999,0,44.15,0,0,Offer B,47758,1,0,0,1,43,0,0.0,0.0,0.0,1931.3,0,1,90247
6684,0,0,0,1,11,0,No phone service,DSL,1,0,0,0,One year,1,Mailed check,36.05,402.6,0,54,17,0.0,4265,0,Gardena,0,0,Cable,33.876482,-118.284077,0,36.05,1,0,None,9960,1,0,0,0,11,1,68.0,0.0,0.0,402.6,0,0,90248
6685,0,0,1,0,45,1,0,DSL,0,0,0,0,Month-to-month,1,Credit card (automatic),50.25,2221.55,0,42,22,6.49,2036,0,Gardena,1,0,Fiber Optic,33.90139,-118.315697,1,50.25,0,6,Offer B,26442,0,0,1,0,45,0,48.87,292.05,0.0,2221.55,0,1,90249
6686,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),109.75,7758.9,0,53,17,22.95,5791,0,Hawthorne,1,1,Fiber Optic,33.914775,-118.348083,1,109.75,0,6,None,93315,1,0,1,1,72,2,1319.0,1652.4,0.0,7758.9,0,0,90250
6687,0,1,1,0,2,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,79.2,172.85,1,78,20,17.73,4225,1,Hermosa Beach,1,0,Cable,33.865320000000004,-118.396336,1,82.36800000000002,0,1,Offer E,18693,0,0,1,0,2,1,35.0,35.46,0.0,172.85,0,0,90254
6688,0,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.3,224.5,0,48,0,19.28,5190,0,Huntington Park,0,0,NA,33.97803,-118.217141,1,20.3,3,3,None,78114,0,0,1,0,12,0,0.0,231.36,0.0,224.5,0,0,90255
6689,0,0,1,1,67,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),112.35,7388.45,0,20,52,20.41,5427,0,Lawndale,1,0,Cable,33.88856,-118.35181299999999,1,112.35,3,3,None,33300,1,0,1,1,67,0,0.0,1367.47,0.0,7388.45,1,1,90260
6690,1,0,1,0,37,1,1,Fiber optic,0,0,1,0,Two year,0,Mailed check,94.3,3460.95,0,23,58,13.13,2615,0,Lynwood,1,1,Fiber Optic,33.923573,-118.20066899999999,1,94.3,0,8,Offer C,69850,1,0,1,0,37,0,0.0,485.81,0.0,3460.95,1,1,90262
6691,0,0,0,0,39,0,No phone service,DSL,1,1,0,0,One year,0,Bank transfer (automatic),41.15,1700.9,0,19,73,0.0,3445,0,Malibu,0,0,DSL,34.037037,-118.705803,0,41.15,0,0,Offer C,11,1,0,0,0,39,0,1242.0,0.0,0.0,1700.9,1,0,90263
6692,0,0,0,0,41,1,1,DSL,1,0,0,1,Month-to-month,1,Bank transfer (automatic),74.65,3090.65,0,47,12,31.08,3859,0,Malibu,1,0,DSL,34.074571999999996,-118.831181,0,74.65,0,0,Offer B,19630,1,0,0,1,41,0,0.0,1274.28,0.0,3090.65,0,1,90265
6693,0,0,0,0,25,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,48.25,1293.8,0,20,59,0.0,4284,0,Manhattan Beach,1,0,DSL,33.889632,-118.39737,0,48.25,0,0,Offer C,33758,0,2,0,1,25,2,763.0,0.0,0.0,1293.8,1,0,90266
6694,1,0,1,1,8,1,1,DSL,1,1,0,1,Two year,1,Credit card (automatic),76.15,645.8,0,32,14,37.28,4457,0,Maywood,0,1,DSL,33.988572,-118.18656499999999,1,76.15,1,0,Offer E,28094,1,0,0,1,8,0,90.0,298.24,0.0,645.8,0,0,90270
6695,0,0,1,1,71,1,1,DSL,1,1,0,0,Two year,0,Mailed check,71.1,5224.95,0,63,52,45.81,6090,0,Pacific Palisades,1,0,DSL,34.079449,-118.54830600000001,1,71.1,3,9,None,22548,1,0,1,0,71,2,2717.0,3252.51,0.0,5224.95,0,0,90272
6696,1,0,0,0,5,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Electronic check,96.55,500.1,0,40,20,39.13,3787,0,Palos Verdes Peninsula,1,1,Cable,33.788208000000004,-118.404955,0,96.55,0,0,None,24979,0,0,0,1,5,0,0.0,195.65,0.0,500.1,0,1,90274
6697,0,0,0,0,30,1,1,DSL,1,0,1,1,One year,1,Credit card (automatic),79.3,2427.1,0,59,18,6.74,2655,0,Rancho Palos Verdes,1,0,Fiber Optic,33.753146,-118.36745900000001,0,79.3,0,0,Offer C,41263,0,0,0,1,30,2,437.0,202.2,0.0,2427.1,0,0,90275
6698,1,0,0,0,40,1,0,Fiber optic,0,1,0,1,One year,1,Credit card (automatic),89.6,3488.15,0,30,69,32.27,2524,0,Redondo Beach,0,1,Cable,33.830453000000006,-118.384565,0,89.6,0,0,Offer B,34191,1,0,0,1,40,0,2407.0,1290.8000000000004,0.0,3488.15,0,0,90277
6699,0,0,0,0,54,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.5,1035.7,0,44,0,10.83,5946,0,Redondo Beach,0,0,NA,33.873395,-118.37019,0,20.5,0,0,Offer B,37322,0,1,0,0,54,1,0.0,584.82,0.0,1035.7,0,0,90278
6700,1,0,1,0,72,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),106.3,7565.35,0,22,85,15.09,4634,0,South Gate,1,1,Fiber Optic,33.944624,-118.19261499999999,1,106.3,0,10,None,96267,0,0,1,1,72,3,6431.0,1086.48,0.0,7565.35,1,0,90280
6701,1,0,1,1,28,1,0,Fiber optic,0,1,1,1,One year,0,Bank transfer (automatic),100.35,2799,0,39,13,7.73,3411,0,Topanga,1,1,DSL,34.115192,-118.61017,1,100.35,2,8,None,5451,0,0,1,1,28,0,364.0,216.44,0.0,2799.0,0,0,90290
6702,1,0,1,1,18,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.6,1601.5,0,45,28,28.04,5968,0,Venice,0,1,Cable,33.991782,-118.479229,1,85.6,3,1,None,31021,1,0,1,1,18,2,0.0,504.72,0.0,1601.5,0,1,90291
6703,0,0,0,0,2,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,45.25,85.5,1,28,53,0.0,4566,1,Marina Del Rey,0,0,Fiber Optic,33.977468,-118.445475,0,47.06,0,0,None,18058,0,4,0,1,2,1,45.0,0.0,0.0,85.5,1,0,90292
6704,0,0,1,1,59,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,106.15,6256.2,0,63,19,35.23,5096,0,Playa Del Rey,1,0,DSL,33.947305,-118.43984099999999,1,106.15,1,1,Offer B,11264,0,0,1,1,59,1,1189.0,2078.57,0.0,6256.2,0,0,90293
6705,1,0,1,1,22,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,51.1,1232.9,0,29,27,27.91,5329,0,Inglewood,0,1,Fiber Optic,33.956445,-118.35863400000001,1,51.1,2,3,None,37527,1,0,1,0,22,0,333.0,614.02,0.0,1232.9,1,0,90301
6706,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.9,19.9,0,55,0,2.38,4050,0,Inglewood,0,0,NA,33.975332,-118.35525200000001,0,19.9,0,0,None,30779,0,0,0,0,1,0,0.0,2.38,0.0,19.9,0,0,90302
6707,0,1,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),25.7,1937.4,0,70,0,8.48,5079,0,Inglewood,0,0,NA,33.936291,-118.33263899999999,1,25.7,0,9,None,27778,0,1,1,0,72,2,0.0,610.5600000000002,0.0,1937.4,0,0,90303
6708,0,1,0,0,14,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.3,1096.25,1,75,11,35.07,5342,1,Inglewood,0,0,DSL,33.936827,-118.359824,0,77.27199999999999,0,0,None,28680,0,1,0,0,14,3,0.0,490.98,0.0,1096.25,0,1,90304
6709,1,0,1,0,50,1,1,Fiber optic,0,0,1,1,One year,0,Electronic check,99.4,5059.75,0,44,18,26.06,6479,0,Inglewood,0,1,Cable,33.958134,-118.330905,1,99.4,0,7,Offer B,13779,1,0,1,1,50,1,0.0,1303.0,0.0,5059.75,0,1,90305
6710,0,0,1,1,48,1,0,DSL,1,0,1,0,One year,0,Bank transfer (automatic),69.7,3023.65,0,19,27,44.66,3442,0,Santa Monica,1,0,Fiber Optic,34.015481,-118.49323100000001,1,69.7,1,6,Offer B,5221,1,0,1,0,48,0,0.0,2143.68,0.0,3023.65,1,1,90401
6711,0,0,1,1,49,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,98.35,4889.2,0,52,57,27.38,4325,0,Santa Monica,0,0,Fiber Optic,34.035849,-118.50350800000001,1,98.35,3,7,Offer B,11509,0,0,1,1,49,2,2787.0,1341.62,0.0,4889.2,0,0,90402
6712,1,0,1,1,28,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,85.45,2289.9,0,64,12,3.18,4022,0,Santa Monica,1,1,Fiber Optic,34.031529,-118.491156,1,85.45,2,6,None,23559,0,0,1,0,28,1,275.0,89.04,0.0,2289.9,0,0,90403
6713,1,1,0,0,68,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,95.9,6503.2,0,66,28,19.67,5080,0,Santa Monica,1,1,Fiber Optic,34.026334000000006,-118.474222,0,95.9,0,0,None,19975,0,0,0,0,68,0,1821.0,1337.5600000000004,0.0,6503.2,0,0,90404
6714,1,0,0,0,13,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,100.75,1313.25,0,29,41,44.43,5985,0,Santa Monica,0,1,Fiber Optic,34.005439,-118.477507,0,100.75,0,0,Offer D,26099,1,0,0,1,13,0,0.0,577.59,0.0,1313.25,1,1,90405
6715,0,0,0,0,11,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,89.2,990.3,0,60,29,10.95,3734,0,Torrance,1,0,Fiber Optic,33.833698999999996,-118.31438700000001,0,89.2,0,0,Offer D,40705,0,0,0,0,11,0,28.72,120.45,0.0,990.3,0,1,90501
6716,0,0,1,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),74.1,228,1,55,26,16.29,5657,1,Torrance,0,0,Cable,33.833181,-118.29206200000002,1,77.064,0,1,None,17058,0,0,1,0,3,5,59.0,48.87,0.0,228.0,0,0,90502
6717,1,1,1,0,57,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,100.6,5746.15,1,73,3,42.1,5247,1,Torrance,1,1,Cable,33.840399,-118.353714,1,104.624,0,1,Offer B,41979,0,3,1,0,57,4,0.0,2399.7000000000007,0.0,5746.15,0,1,90503
6718,1,0,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Mailed check,75.0,209.1,1,27,57,34.49,3190,1,Torrance,0,1,Cable,33.867257,-118.330794,0,78.0,0,0,None,31678,0,0,0,1,3,3,119.0,103.47,0.0,209.1,1,0,90504
6719,1,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.75,1864.2,0,62,0,40.04,4413,0,Torrance,0,1,NA,33.807882,-118.34795700000001,1,25.75,0,1,None,34873,0,0,1,0,72,0,0.0,2882.88,0.0,1864.2,0,0,90505
6720,1,0,1,1,70,1,1,DSL,0,1,1,1,Two year,1,Electronic check,84.1,5979.7,0,63,24,38.83,5568,0,Whittier,1,1,DSL,34.007353,-118.03368300000001,1,84.1,3,4,None,32050,1,0,1,1,70,2,1435.0,2718.1,0.0,5979.7,0,0,90601
6721,0,0,1,1,49,1,1,DSL,0,1,1,1,Two year,0,Bank transfer (automatic),79.3,3902.45,0,47,14,16.6,6366,0,Whittier,0,0,Fiber Optic,33.972119,-118.02018799999999,1,79.3,1,9,Offer B,26265,1,2,1,1,49,2,546.0,813.4000000000002,0.0,3902.45,0,0,90602
6722,0,1,1,0,67,1,1,Fiber optic,1,0,1,1,One year,1,Credit card (automatic),107.05,7142.5,0,67,20,38.47,4126,0,Whittier,1,0,Fiber Optic,33.945318,-117.992066,1,107.05,0,8,None,19109,0,0,1,0,67,1,0.0,2577.49,0.0,7142.5,0,1,90603
6723,1,0,0,0,46,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.05,902,0,61,0,30.25,2942,0,Whittier,0,1,NA,33.929704,-118.01208000000001,0,20.05,0,0,Offer B,37887,0,0,0,0,46,0,0.0,1391.5,0.0,902.0,0,0,90604
6724,0,1,0,0,64,1,0,DSL,1,1,1,0,Two year,1,Credit card (automatic),70.2,4481,1,80,26,29.12,6080,1,Whittier,0,0,Cable,33.960891,-118.03222199999999,0,73.00800000000002,0,0,Offer B,38181,1,0,0,0,64,1,1165.0,1863.68,0.0,4481.0,0,0,90605
6725,0,0,1,0,37,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),19.5,805.2,0,57,0,45.19,3924,0,Whittier,0,0,NA,33.976678,-118.065875,1,19.5,0,1,None,32148,0,0,1,0,37,2,0.0,1672.03,0.0,805.2,0,0,90606
6726,0,1,0,0,2,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,70.75,154.85,1,74,23,9.86,4407,1,Buena Park,0,0,Cable,33.845706,-118.012204,0,73.58,0,0,Offer E,44442,0,0,0,0,2,3,36.0,19.72,0.0,154.85,0,0,90620
6727,0,1,1,0,13,0,No phone service,DSL,0,0,1,1,Month-to-month,0,Electronic check,45.3,528.45,0,68,9,0.0,4118,0,Buena Park,0,0,Fiber Optic,33.874224,-117.99336799999999,1,45.3,0,5,None,33528,0,0,1,0,13,0,4.76,0.0,0.0,528.45,0,1,90621
6728,0,0,1,0,72,1,1,Fiber optic,1,1,1,1,Two year,0,Electronic check,115.15,8349.7,0,63,25,40.59,4761,0,La Palma,1,0,DSL,33.850504,-118.039892,1,115.15,0,10,None,15505,1,0,1,1,72,0,0.0,2922.4800000000005,0.0,8349.7,0,1,90623
6729,1,0,1,1,68,1,0,DSL,0,0,1,1,Two year,1,Bank transfer (automatic),72.95,4953.25,0,45,25,34.13,4499,0,Cypress,1,1,DSL,33.818477,-118.038307,1,72.95,1,4,None,47344,1,2,1,1,68,1,0.0,2320.84,0.0,4953.25,0,1,90630
6730,1,0,1,1,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.65,332.65,0,48,0,17.28,5928,0,La Habra,0,1,NA,33.940619,-117.9513,1,19.65,3,1,Offer D,67354,0,0,1,0,15,0,0.0,259.20000000000005,0.0,332.65,0,0,90631
6731,0,0,0,0,24,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.55,470.2,0,51,0,10.64,2511,0,La Mirada,0,0,NA,33.902045,-118.00896100000001,0,19.55,0,0,None,47568,0,1,0,0,24,3,0.0,255.36,0.0,470.2,0,0,90638
6732,0,0,0,0,24,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.55,2259.35,0,21,52,18.07,5352,0,Montebello,0,0,Cable,34.015217,-118.10996200000001,0,89.55,0,0,None,62425,1,0,0,1,24,0,0.0,433.68,0.0,2259.35,1,1,90640
6733,1,0,0,0,27,1,0,DSL,1,0,0,0,Month-to-month,0,Mailed check,50.35,1411.35,0,59,9,18.51,5578,0,Norwalk,0,1,Fiber Optic,33.905963,-118.08263000000001,0,50.35,0,0,None,103214,0,0,0,0,27,3,0.0,499.77,0.0,1411.35,0,1,90650
6734,1,0,0,0,12,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),50.25,593.75,1,50,29,46.58,3624,1,Pico Rivera,0,1,Fiber Optic,33.989523999999996,-118.089299,0,52.26000000000001,0,0,None,63288,1,0,0,0,12,1,0.0,558.96,0.0,593.75,0,1,90660
6735,0,0,1,1,71,1,0,DSL,1,1,1,1,Two year,0,Credit card (automatic),87.25,6328.7,0,24,51,48.08,4135,0,Santa Fe Springs,1,0,DSL,33.933565,-118.062611,1,87.25,2,5,None,16271,1,0,1,1,71,2,322.76,3413.68,0.0,6328.7,1,1,90670
6736,1,0,1,1,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.8,1411.9,0,48,0,8.82,5626,0,Stanton,0,1,NA,33.801869,-117.99506799999999,1,20.8,2,6,None,29694,0,0,1,0,67,0,0.0,590.94,0.0,1411.9,0,0,90680
6737,0,0,1,0,63,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),109.25,6841.4,0,64,23,10.67,5700,0,Artesia,1,0,DSL,33.867593,-118.08063700000001,1,109.25,0,8,None,16398,1,2,1,1,63,2,157.35,672.21,0.0,6841.4,0,1,90701
6738,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.35,20.35,0,50,0,31.97,2648,0,Cerritos,0,1,NA,33.8681,-118.067402,0,20.35,0,0,None,51556,0,0,0,0,1,1,0.0,31.97,0.0,20.35,0,0,90703
6739,1,0,0,0,4,1,0,DSL,0,0,0,1,Month-to-month,1,Electronic check,55.9,238.5,0,51,22,17.7,3545,0,Avalon,0,1,DSL,33.391181,-118.421305,0,55.9,0,0,None,3699,0,0,0,1,4,2,52.0,70.8,0.0,238.5,0,0,90704
6740,0,1,0,0,40,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),79.2,3233.85,1,65,4,44.86,3207,1,Bellflower,0,0,Fiber Optic,33.887676,-118.12728899999999,0,82.36800000000002,0,0,Offer B,72893,0,0,0,0,40,3,0.0,1794.4,0.0,3233.85,0,1,90706
6741,0,0,0,0,12,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,96.0,1062.1,1,46,30,25.54,5239,1,Harbor City,1,0,Fiber Optic,33.798266,-118.30023700000001,0,99.84,0,0,None,24660,0,0,0,1,12,0,0.0,306.48,0.0,1062.1,0,1,90710
6742,1,0,1,1,52,1,0,DSL,1,1,1,1,Two year,0,Electronic check,79.2,4016.3,0,61,12,16.53,4509,0,Lakewood,1,1,Fiber Optic,33.840524,-118.148403,1,79.2,2,5,None,30173,0,0,1,1,52,0,0.0,859.5600000000002,0.0,4016.3,0,1,90712
6743,1,0,0,0,10,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,24.0,226.55,0,35,0,3.01,5299,0,Lakewood,0,1,NA,33.847755,-118.112532,0,24.0,0,0,Offer D,27563,0,1,0,0,10,3,0.0,30.1,0.0,226.55,0,0,90713
6744,1,0,0,0,68,1,1,Fiber optic,1,1,1,0,One year,0,Bank transfer (automatic),101.35,7110.75,0,56,7,11.22,4941,0,Lakewood,1,1,Cable,33.841027000000004,-118.078097,0,101.35,0,0,None,20890,0,0,0,0,68,0,498.0,762.96,0.0,7110.75,0,0,90715
6745,0,0,0,0,54,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.1,5440.9,1,38,10,41.83,5763,1,Hawaiian Gardens,0,0,Fiber Optic,33.830431,-118.07407099999999,0,104.104,0,0,None,14852,1,3,0,1,54,2,0.0,2258.82,0.0,5440.9,0,1,90716
6746,0,0,1,1,4,1,0,DSL,0,1,0,0,Month-to-month,0,Mailed check,56.5,235.1,1,38,62,42.71,5758,1,Lomita,0,0,DSL,33.794209,-118.31735400000001,1,58.76000000000001,3,5,None,21065,1,0,1,0,4,4,0.0,170.84,0.0,235.1,0,1,90717
6747,0,0,1,0,52,0,No phone service,DSL,1,0,0,0,One year,0,Mailed check,35.45,1958.95,0,58,8,0.0,5509,0,Los Alamitos,1,0,Fiber Optic,33.794990000000006,-118.065591,1,35.45,0,4,None,21343,0,0,1,0,52,1,157.0,0.0,0.0,1958.95,0,0,90720
6748,0,1,0,0,1,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,85.0,85,1,71,9,42.5,2650,1,Paramount,1,0,Cable,33.897121999999996,-118.164432,0,88.4,0,0,None,55306,0,2,0,0,1,2,0.0,42.5,0.0,85.0,0,0,90723
6749,1,0,1,0,70,1,1,DSL,1,1,1,0,One year,0,Bank transfer (automatic),79.4,5528.9,0,40,21,43.46,5991,0,San Pedro,1,1,Fiber Optic,33.736387,-118.28436299999998,1,79.4,0,0,None,58639,1,1,0,0,70,1,0.0,3042.2000000000007,0.0,5528.9,0,1,90731
6750,1,0,0,0,43,0,No phone service,DSL,1,0,0,0,One year,1,Credit card (automatic),35.2,1463.7,0,47,4,0.0,5268,0,San Pedro,1,1,Fiber Optic,33.744119,-118.31448,0,35.2,0,0,None,21279,0,0,0,0,43,1,59.0,0.0,0.0,1463.7,0,0,90732
6751,1,0,0,0,52,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.65,1025.05,0,31,0,21.98,5157,0,Seal Beach,0,1,NA,33.75462,-118.071128,0,19.65,0,0,None,24180,0,0,0,0,52,0,0.0,1142.96,0.0,1025.05,0,0,90740
6752,0,0,0,0,12,0,No phone service,DSL,1,0,0,1,Two year,0,Mailed check,49.85,552.1,0,58,7,0.0,3100,0,Sunset Beach,1,0,Cable,33.719221000000005,-118.073596,0,49.85,0,0,Offer D,1107,1,0,0,1,12,0,0.0,0.0,0.0,552.1,0,1,90742
6753,0,0,1,1,56,1,1,DSL,1,1,0,1,One year,0,Bank transfer (automatic),68.75,3815.4,0,25,76,7.31,6494,0,Surfside,0,0,Fiber Optic,33.728273,-118.08530400000001,1,68.75,1,7,None,174,0,0,1,1,56,0,0.0,409.36,0.0,3815.4,1,1,90743
6754,1,0,0,1,0,1,1,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),61.9, ,0,56,19,29.95,5188,0,Wilmington,0,1,Cable,33.782068,-118.26226299999999,0,61.9,1,0,None,53323,1,0,0,0,10,0,0.0,299.5,0.0,619.0,0,1,90744
6755,1,0,0,0,42,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,79.9,3313.4,0,53,14,9.46,2583,0,Carson,1,1,DSL,33.822295000000004,-118.26411,0,79.9,0,0,None,55486,0,0,0,0,42,1,46.39,397.32000000000005,23.47,3313.4,0,1,90745
6756,1,1,1,0,22,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),89.75,1938.9,0,65,14,22.38,4180,0,Carson,0,1,Fiber Optic,33.859171,-118.25227199999999,1,89.75,0,8,None,25566,0,0,1,1,22,0,0.0,492.36,0.0,1938.9,0,1,90746
6757,1,0,1,1,51,0,No phone service,DSL,1,1,1,1,One year,0,Electronic check,59.3,3014.65,1,51,2,0.0,5633,1,Long Beach,1,1,Fiber Optic,33.752524,-118.21073700000001,1,61.672,0,1,None,38427,0,0,1,1,51,2,60.0,0.0,0.0,3014.65,0,0,90802
6758,1,0,0,0,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),19.4,460.25,0,43,0,2.59,5975,0,Long Beach,0,1,NA,33.760458,-118.129725,0,19.4,0,0,None,31352,0,0,0,0,27,1,0.0,69.92999999999999,29.59,460.25,0,0,90803
6759,1,1,1,0,51,1,1,Fiber optic,1,0,0,1,One year,1,Bank transfer (automatic),93.65,4839.15,0,76,10,2.21,4163,0,Long Beach,1,1,Fiber Optic,33.783046999999996,-118.1486,1,93.65,0,7,Offer B,43467,0,0,1,0,51,2,484.0,112.71,0.0,4839.15,0,0,90804
6760,1,0,0,1,4,1,0,DSL,1,0,0,0,Month-to-month,1,Electronic check,49.4,184.4,1,44,18,9.77,4455,1,Long Beach,0,1,DSL,33.864622,-118.179626,0,51.376000000000005,2,0,None,91664,0,0,0,0,4,4,33.0,39.08,0.0,184.4,0,0,90805
6761,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.9,19.9,0,36,0,7.76,4590,0,Long Beach,0,1,NA,33.802664,-118.179971,0,19.9,0,0,None,49647,0,1,0,0,1,2,0.0,7.76,0.0,19.9,0,0,90806
6762,1,0,0,0,35,1,0,DSL,0,0,1,0,Month-to-month,0,Mailed check,55.0,2010.55,1,60,15,48.93,2220,1,Long Beach,0,1,Cable,33.830099,-118.182239,0,57.2,0,0,None,31556,0,0,0,0,35,2,302.0,1712.55,0.0,2010.55,0,0,90807
6763,1,1,1,1,71,1,1,DSL,0,1,0,1,One year,1,Bank transfer (automatic),72.9,5139.65,0,74,20,46.11,6404,0,Long Beach,1,1,Fiber Optic,33.823943,-118.11133500000001,1,72.9,3,1,None,37417,1,1,1,0,71,1,1028.0,3273.81,0.0,5139.65,0,0,90808
6764,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.2,69.2,1,51,20,10.08,2637,1,Long Beach,0,0,Fiber Optic,33.819814,-118.222416,0,71.968,0,0,None,35656,0,0,0,0,1,6,0.0,10.08,0.0,69.2,0,0,90810
6765,0,0,1,1,69,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.6,1673.4,0,55,0,20.98,6053,0,Long Beach,0,0,NA,33.781086,-118.199049,1,25.6,1,5,None,63136,0,0,1,0,69,0,0.0,1447.62,28.09,1673.4,0,0,90813
6766,1,0,1,1,14,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,19.75,309.35,0,38,0,26.99,3958,0,Long Beach,0,1,NA,33.771612,-118.14386599999999,1,19.75,2,6,Offer D,19034,0,0,1,0,14,0,0.0,377.86,6.49,309.35,0,0,90814
6767,1,0,1,0,57,1,0,DSL,1,0,0,0,Month-to-month,0,Electronic check,55.7,3171.6,0,31,15,15.48,4607,0,Long Beach,0,1,DSL,33.797638,-118.11662,1,55.7,0,6,None,38902,1,0,1,0,57,2,476.0,882.36,34.59,3171.6,0,0,90815
6768,0,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,0,Credit card (automatic),117.5,8670.1,0,58,16,33.37,6009,0,Long Beach,1,0,Fiber Optic,33.778436,-118.118648,1,117.5,1,9,None,425,1,0,1,1,72,3,1387.0,2402.64,47.55,8670.1,0,0,90822
6769,1,0,0,0,48,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.85,916,0,63,0,32.04,3779,0,Altadena,0,1,NA,34.196837,-118.14223600000001,0,19.85,0,0,None,36243,0,0,0,0,48,2,0.0,1537.92,0.0,916.0,0,0,91001
6770,0,0,1,1,4,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,78.9,299.75,0,35,53,41.93,5775,0,Arcadia,0,0,Cable,34.137319,-118.02983700000001,1,78.9,3,9,None,30028,0,2,1,0,4,2,0.0,167.72,37.01,299.75,0,1,91006
6771,1,0,1,1,31,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,20.65,702.05,0,31,0,9.56,2990,0,Arcadia,0,1,NA,34.128284,-118.04773200000001,1,20.65,1,10,None,30933,0,0,1,0,31,1,0.0,296.36,43.76,702.05,0,0,91007
6772,1,0,0,0,38,1,0,DSL,0,0,0,1,One year,1,Mailed check,62.3,2354.8,1,46,15,46.21,3818,1,Duarte,1,1,Cable,34.145695,-117.95982,0,64.792,0,0,None,27414,1,0,0,1,38,2,353.0,1755.98,0.0,2354.8,0,0,91010
6773,1,1,1,0,37,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,92.5,3473.4,1,74,4,49.37,4127,1,La Canada Flintridge,0,1,Cable,34.234912,-118.153729,1,96.2,0,3,None,20200,0,3,1,1,37,1,0.0,1826.69,0.0,3473.4,0,1,91011
6774,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,19.65,19.65,0,28,0,42.42,5454,0,Monrovia,0,0,NA,34.1528,-118.000482,0,19.65,0,0,None,41067,0,0,0,0,1,0,0.0,42.42,0.0,19.65,1,0,91016
6775,1,1,0,0,57,1,1,DSL,0,1,1,1,Two year,1,Bank transfer (automatic),79.75,4438.2,0,72,16,9.1,5371,0,Montrose,1,1,Cable,34.2112,-118.230625,0,79.75,0,0,Offer B,7527,0,0,0,0,57,2,710.0,518.6999999999998,0.0,4438.2,0,0,91020
6776,0,1,1,0,62,1,0,DSL,1,0,1,1,Two year,1,Credit card (automatic),79.95,4819.75,0,69,29,24.62,6488,0,Sierra Madre,1,0,Cable,34.168686,-118.057505,1,79.95,0,9,Offer B,10558,1,0,1,0,62,2,0.0,1526.44,0.0,4819.75,0,1,91024
6777,1,0,1,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,29.9,92.25,0,22,41,0.0,4416,0,South Pasadena,0,1,Fiber Optic,34.110444,-118.156957,1,29.9,0,5,None,23984,1,0,1,0,3,1,38.0,0.0,0.0,92.25,1,0,91030
6778,0,0,0,1,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,19.75,1567,0,56,0,15.21,5478,0,Sunland,0,0,NA,34.282703999999995,-118.312929,0,19.75,2,0,None,18752,0,0,0,0,72,1,0.0,1095.12,25.98,1567.0,0,0,91040
6779,1,0,0,1,29,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Mailed check,45.0,1242.45,0,57,21,0.0,3290,0,Tujunga,1,1,DSL,34.296574,-118.24483899999998,0,45.0,1,0,None,26753,1,0,0,0,29,0,261.0,0.0,12.26,1242.45,0,0,91042
6780,1,0,1,1,13,1,0,DSL,0,0,0,0,Month-to-month,0,Bank transfer (automatic),44.8,559.2,0,25,59,6.18,4680,0,Pasadena,0,1,DSL,34.146634999999996,-118.139225,1,44.8,3,0,None,16812,0,0,0,0,13,0,32.99,80.34,37.49,559.2,1,1,91101
6781,1,0,0,1,3,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,69.65,220.1,1,53,25,39.38,2421,1,Pasadena,0,1,Fiber Optic,34.167465,-118.165327,0,72.436,0,0,Offer E,27891,0,0,0,0,3,0,55.0,118.14,0.0,220.1,0,0,91103
6782,0,0,0,0,11,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,51.1,531.15,0,64,21,2.95,4467,0,Pasadena,0,0,DSL,34.165383,-118.123752,0,51.1,0,0,None,38460,0,0,0,0,11,1,0.0,32.45,0.0,531.15,0,1,91104
6783,0,0,0,1,21,0,No phone service,DSL,1,1,1,0,Two year,0,Mailed check,53.15,1183.2,0,59,11,0.0,3461,0,Pasadena,1,0,Fiber Optic,34.13946,-118.16664899999999,0,53.15,1,0,None,10253,1,0,0,0,21,3,0.0,0.0,19.13,1183.2,0,1,91105
6784,0,0,0,0,19,1,1,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Bank transfer (automatic),24.7,465.85,0,62,0,11.86,3612,0,Pasadena,0,0,NA,34.139402000000004,-118.128658,0,24.7,0,0,None,23742,0,0,0,0,19,0,0.0,225.34,1.65,465.85,0,0,91106
6785,1,0,0,0,61,1,1,Fiber optic,1,0,1,1,Two year,1,Credit card (automatic),111.6,6876.05,1,44,12,7.82,4495,1,Pasadena,1,1,DSL,34.159007,-118.08735300000001,0,116.064,0,0,None,32369,1,1,0,1,61,2,0.0,477.02,0.0,6876.05,0,1,91107
6786,0,0,0,0,11,1,0,DSL,1,0,0,0,Month-to-month,0,Credit card (automatic),48.55,501,1,43,9,19.01,4444,1,San Marino,0,0,Cable,34.122671000000004,-118.11291100000001,0,50.492,0,0,None,13158,0,0,0,0,11,2,0.0,209.11,0.0,501.0,0,1,91108
6787,1,0,1,1,35,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,109.95,3782.4,0,24,73,48.3,5721,0,Glendale,1,1,DSL,34.17051,-118.28946299999998,1,109.95,3,8,None,23981,1,0,1,1,35,0,0.0,1690.5,31.9,3782.4,1,1,91201
6788,1,0,0,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.8,460.2,0,55,0,3.07,3274,0,Glendale,0,1,NA,34.167926,-118.26753899999999,0,20.8,3,0,None,21990,0,0,0,0,25,0,0.0,76.75,21.81,460.2,0,0,91202
6789,0,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.2,20.2,1,62,0,48.25,4197,1,Glendale,0,0,NA,34.153338,-118.262974,0,20.2,0,0,Offer E,14493,0,0,0,0,1,3,0.0,48.25,0.0,20.2,0,0,91203
6790,0,0,0,0,67,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),25.6,1790.35,0,53,0,16.72,5183,0,Glendale,0,0,NA,34.136306,-118.26036,0,25.6,0,0,None,17015,0,0,0,0,67,1,0.0,1120.24,46.06,1790.35,0,0,91204
6791,1,0,0,0,19,0,No phone service,DSL,0,0,1,0,Month-to-month,1,Electronic check,39.65,733.35,1,50,23,0.0,2933,1,Glendale,1,1,Fiber Optic,34.13658,-118.24583899999999,0,41.236000000000004,0,0,None,41390,0,3,0,0,19,6,169.0,0.0,0.0,733.35,0,0,91205
6792,1,0,0,0,56,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,24.9,1334,1,57,0,2.58,5327,1,Glendale,0,1,NA,34.162515,-118.203869,0,24.9,0,0,None,31297,0,0,0,0,56,2,0.0,144.48000000000005,0.0,1334.0,0,0,91206
6793,1,0,1,1,72,1,1,Fiber optic,1,1,1,1,Two year,1,Credit card (automatic),108.4,7767.25,0,56,30,27.88,4419,0,Glendale,1,1,Fiber Optic,34.182378,-118.262922,1,108.4,2,4,None,9864,0,0,1,1,72,1,0.0,2007.36,0.0,7767.25,0,1,91207
6794,1,0,0,0,43,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.55,876.15,0,57,0,3.18,4871,0,Glendale,0,1,NA,34.195386,-118.23850800000001,0,19.55,0,0,None,16910,0,0,0,0,43,0,0.0,136.74,15.17,876.15,0,0,91208
6795,0,0,1,1,55,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Electronic check,85.1,4600.95,0,51,19,20.1,4026,0,La Crescenta,0,0,Fiber Optic,34.239636,-118.245259,1,85.1,2,5,None,29110,0,0,1,0,55,1,874.0,1105.5,14.3,4600.95,0,0,91214
6796,1,0,1,1,2,1,1,DSL,1,0,0,0,Month-to-month,0,Mailed check,56.7,113.55,1,62,58,5.67,5560,1,Agoura Hills,0,1,Cable,34.129058,-118.75978799999999,1,58.968,3,1,None,25303,0,0,1,0,2,2,0.0,11.34,0.0,113.55,0,1,91301
6797,1,0,0,0,27,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,69.05,1793.25,0,26,26,34.98,3241,0,Calabasas,0,1,Cable,34.130860999999996,-118.68346000000001,0,69.05,0,0,None,23661,0,0,0,0,27,0,466.0,944.46,22.72,1793.25,1,0,91302
6798,0,0,0,0,13,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.15,886.7,0,40,28,26.13,2992,0,Canoga Park,0,0,Fiber Optic,34.19829,-118.602203,0,70.15,0,0,None,23519,0,0,0,0,13,2,248.0,339.69,8.53,886.7,0,0,91303
6799,0,0,0,0,70,1,1,Fiber optic,1,1,1,1,Two year,1,Mailed check,111.15,7737.55,0,63,17,23.15,4240,0,Canoga Park,1,0,Fiber Optic,34.224377000000004,-118.63265600000001,0,111.15,0,0,None,49242,0,0,0,1,70,0,1315.0,1620.5,46.26,7737.55,0,0,91304
6800,0,0,1,0,14,1,0,Fiber optic,1,1,1,1,One year,0,Mailed check,105.95,1348.9,1,59,25,5.63,5887,1,Winnetka,0,0,Cable,34.209532,-118.57756299999998,1,110.18799999999999,0,3,None,43857,1,0,1,1,14,4,0.0,78.82,0.0,1348.9,0,1,91306
6801,0,0,1,1,19,1,1,Fiber optic,0,0,0,1,One year,1,Bank transfer (automatic),89.35,1686.85,0,24,52,36.92,4473,0,West Hills,0,0,Fiber Optic,34.199787,-118.68493000000001,1,89.35,3,1,None,23637,1,2,1,1,19,1,0.0,701.48,0.0,1686.85,1,1,91307
6802,0,0,0,0,20,1,1,Fiber optic,1,0,1,0,Month-to-month,1,Bank transfer (automatic),89.1,1879.25,0,50,25,24.73,3027,0,Chatsworth,0,0,Fiber Optic,34.294142,-118.60388300000001,0,89.1,0,0,None,35325,0,0,0,0,20,0,46.98,494.6,15.43,1879.25,0,1,91311
6803,1,0,1,1,43,1,1,Fiber optic,1,0,0,0,One year,1,Credit card (automatic),91.25,4013.8,0,59,25,42.22,5884,0,Encino,1,1,Fiber Optic,34.150354,-118.51829199999999,1,91.25,1,11,None,27614,1,0,1,0,43,2,1003.0,1815.46,25.49,4013.8,0,0,91316
6804,1,0,1,1,5,1,0,Fiber optic,1,0,0,1,Month-to-month,1,Mailed check,90.35,434.5,0,33,19,15.01,4014,0,Newbury Park,1,1,DSL,34.172071,-118.946262,1,90.35,1,1,None,37779,0,1,1,1,5,1,83.0,75.05,17.33,434.5,0,0,91320
6805,0,1,1,0,70,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),105.55,7195.35,0,72,24,33.74,4605,0,Newhall,0,0,Fiber Optic,34.370378,-118.50411799999999,1,105.55,0,1,None,30742,1,0,1,0,70,1,0.0,2361.8,0.0,7195.35,0,1,91321
6806,0,0,1,0,40,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.1,780.1,0,39,0,31.37,2056,0,Northridge,0,0,NA,34.238208,-118.55028999999999,1,19.1,0,1,None,25751,0,0,1,0,40,2,0.0,1254.8,45.6,780.1,0,0,91324
6807,1,0,1,1,6,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.4,107.6,0,54,0,41.36,4628,0,Northridge,0,1,NA,34.236683,-118.51758799999999,1,20.4,3,1,None,32307,0,0,1,0,6,2,0.0,248.16,0.0,107.6,0,0,91325
6808,1,0,0,0,39,1,0,Fiber optic,1,0,1,1,Two year,1,Electronic check,100.45,3801.7,0,38,19,37.94,2698,0,Porter Ranch,1,1,Cable,34.281911,-118.55621799999999,0,100.45,0,0,None,28067,0,0,0,1,39,2,0.0,1479.66,0.0,3801.7,0,1,91326
6809,1,1,1,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,0,Electronic check,74.95,308.7,1,76,30,28.11,3716,1,Pacoima,0,1,DSL,34.255441999999995,-118.421314,1,77.94800000000002,0,1,None,97318,0,0,1,0,4,1,9.26,112.44,0.0,308.7,0,1,91331
6810,1,0,0,0,15,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Electronic check,29.7,438.25,1,56,32,0.0,5518,1,Reseda,0,1,DSL,34.200175,-118.540958,0,30.888,0,0,None,68018,1,0,0,0,15,0,140.0,0.0,0.0,438.25,0,0,91335
6811,1,0,1,0,1,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,50.35,50.35,1,40,22,0.0,4526,1,San Fernando,1,1,DSL,34.286131,-118.435969,1,52.364,0,1,Offer E,33389,0,0,1,1,1,4,0.0,0.0,0.0,50.35,0,0,91340
6812,0,1,0,0,45,1,0,Fiber optic,1,1,0,0,Month-to-month,1,Bank transfer (automatic),85.7,3778.1,0,80,20,4.14,5397,0,Sylmar,0,0,DSL,34.321621,-118.399841,0,85.7,0,0,None,81986,1,0,0,0,45,1,75.56,186.3,0.0,3778.1,0,1,91342
6813,0,0,1,0,64,0,No phone service,DSL,1,0,0,1,Two year,0,Electronic check,47.85,3147.5,1,61,30,0.0,6347,1,North Hills,1,0,DSL,34.238802,-118.48229599999999,1,49.763999999999996,0,5,None,57017,1,0,1,1,64,1,944.0,0.0,0.0,3147.5,0,0,91343
6814,0,1,1,0,57,1,1,Fiber optic,0,1,0,1,Month-to-month,0,Credit card (automatic),94.0,5438.95,0,77,30,23.05,6015,0,Granada Hills,1,0,Fiber Optic,34.291273,-118.505104,1,94.0,0,1,None,48867,0,1,1,0,57,2,0.0,1313.85,0.0,5438.95,0,1,91344
6815,1,0,1,1,72,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),69.85,5102.35,0,62,18,28.37,6233,0,Mission Hills,1,1,DSL,34.266389000000004,-118.459744,1,69.85,2,1,None,17112,1,0,1,0,72,1,0.0,2042.64,25.24,5102.35,0,1,91345
6816,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,70.3,70.3,1,32,8,5.67,4512,1,Santa Clarita,0,1,Fiber Optic,34.502432,-118.41458999999999,0,73.112,0,0,Offer E,40077,0,0,0,0,1,1,0.0,5.67,0.0,70.3,0,0,91350
6817,1,0,1,0,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.85,1872.2,0,36,0,36.03,5514,0,Canyon Country,0,1,NA,34.422519,-118.420717,1,25.85,0,1,None,59259,0,0,1,0,72,4,0.0,2594.16,5.73,1872.2,0,0,91351
6818,0,0,0,0,3,1,0,DSL,1,1,0,1,Two year,0,Mailed check,71.1,213.35,0,36,22,37.0,3501,0,Sun Valley,0,0,Fiber Optic,34.231053,-118.338307,0,71.1,0,0,None,46639,1,0,0,1,3,0,0.0,111.0,2.62,213.35,0,1,91352
6819,1,1,0,0,55,1,1,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,98.8,5617.75,1,73,23,8.93,5543,1,Valencia,0,1,DSL,34.457005,-118.57372600000001,0,102.75200000000001,0,0,Offer B,17846,0,0,0,1,55,1,1292.0,491.15,0.0,5617.75,0,0,91354
6820,0,0,1,0,59,1,1,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,93.35,5386.5,0,45,26,20.78,4814,0,Valencia,1,0,Fiber Optic,34.43987,-118.644609,1,93.35,0,1,None,24977,1,0,1,0,59,0,0.0,1226.02,36.07,5386.5,0,1,91355
6821,0,0,0,0,18,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Bank transfer (automatic),99.85,1776.95,1,34,3,36.49,3068,1,Tarzana,0,0,Fiber Optic,34.157137,-118.548511,0,103.844,0,0,None,27424,1,1,0,1,18,3,0.0,656.82,0.0,1776.95,0,1,91356
6822,1,1,1,0,32,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Credit card (automatic),80.3,2483.05,1,71,28,2.08,5365,1,Thousand Oaks,0,1,Fiber Optic,34.214054,-118.88108999999999,1,83.512,0,1,None,42526,0,1,1,1,32,1,69.53,66.56,0.0,2483.05,0,1,91360
6823,0,0,0,0,4,1,0,DSL,1,0,0,0,Month-to-month,1,Bank transfer (automatic),50.55,235.65,0,24,41,22.07,4164,0,Westlake Village,0,0,DSL,34.130992,-118.894673,0,50.55,0,0,None,18735,0,0,0,0,4,1,97.0,88.28,0.0,235.65,1,0,91361
6824,0,1,0,0,66,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Credit card (automatic),80.45,5224.35,1,72,26,45.59,5011,1,Thousand Oaks,0,0,DSL,34.191842,-118.822796,0,83.66799999999999,0,0,None,33057,0,1,0,0,66,7,1358.0,3008.94,0.0,5224.35,0,0,91362
6825,1,0,0,0,27,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,81.3,2272.8,0,20,69,25.51,5158,0,Woodland Hills,1,1,Cable,34.153733,-118.59340800000001,0,81.3,0,0,None,25988,0,0,0,0,27,2,0.0,688.7700000000002,29.93,2272.8,1,1,91364
6826,1,0,0,0,4,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Credit card (automatic),20.7,83.75,0,49,0,27.04,3027,0,Woodland Hills,0,1,NA,34.178067999999996,-118.61571399999998,0,20.7,0,0,None,36123,0,1,0,0,4,1,0.0,108.16,0.0,83.75,0,0,91367
6827,1,0,1,1,60,1,0,DSL,1,1,1,1,Month-to-month,1,Credit card (automatic),79.05,4663.4,0,59,76,39.76,5275,0,Oak Park,0,1,Cable,34.19225,-118.77687399999999,1,79.05,3,1,None,14814,1,0,1,1,60,0,0.0,2385.6,0.0,4663.4,0,1,91377
6828,0,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,19.05,201.7,0,26,0,42.67,3153,0,Stevenson Ranch,0,0,NA,34.364153,-118.615583,1,19.05,1,1,None,9937,0,1,1,0,8,2,0.0,341.36,0.0,201.7,1,0,91381
6829,1,0,1,1,8,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.6,125,0,54,0,13.43,3214,0,Castaic,0,1,NA,34.506627,-118.699048,1,19.6,3,1,Offer E,22177,0,0,1,0,8,0,0.0,107.44,0.0,125.0,0,0,91384
6830,1,0,0,0,35,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,20.2,684.4,0,64,0,42.8,3481,0,Van Nuys,0,1,NA,34.178483,-118.43179099999999,0,20.2,0,0,None,40376,0,0,0,0,35,3,0.0,1498.0,0.0,684.4,0,0,91401
6831,1,0,0,0,7,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,86.8,620.35,1,22,65,30.61,3780,1,Fallbrook,0,1,Cable,33.362575,-117.299644,0,90.272,0,0,Offer E,42239,0,1,0,1,7,1,403.0,214.27,0.0,620.35,1,0,92028
6832,0,0,1,1,53,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.9,1146.05,0,48,0,43.71,4254,0,Sherman Oaks,0,0,NA,34.147149,-118.463365,1,20.9,3,1,None,22085,0,0,1,0,53,3,0.0,2316.63,0.0,1146.05,0,0,91403
6833,0,1,0,0,18,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),103.6,1806.35,0,65,3,1.27,2094,0,Van Nuys,0,0,Fiber Optic,34.202494,-118.448048,0,103.6,0,0,None,51348,1,0,0,1,18,0,0.0,22.86,0.0,1806.35,0,1,91405
6834,0,0,0,0,15,0,No phone service,DSL,0,1,0,1,Two year,1,Mailed check,38.8,603,0,49,23,0.0,2118,0,Van Nuys,0,0,DSL,34.195685,-118.490752,0,38.8,0,0,None,50047,0,0,0,1,15,1,0.0,0.0,0.0,603.0,0,1,91406
6835,1,0,1,0,67,1,1,Fiber optic,0,1,1,0,One year,1,Bank transfer (automatic),88.4,5798.3,0,44,23,37.6,6251,0,Van Nuys,0,1,Fiber Optic,34.178470000000004,-118.45947199999999,1,88.4,0,1,None,23646,0,1,1,0,67,3,1334.0,2519.2000000000007,0.0,5798.3,0,0,91411
6836,1,1,1,0,6,1,0,Fiber optic,0,1,0,1,Month-to-month,1,Electronic check,84.2,519.15,1,76,28,40.44,5834,1,Sherman Oaks,0,1,Fiber Optic,34.146957,-118.432138,1,87.56800000000001,0,1,None,29387,0,1,1,0,6,2,145.0,242.64,0.0,519.15,0,0,91423
6837,1,1,0,0,6,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,79.7,497.6,0,69,11,48.32,2893,0,Encino,0,1,Fiber Optic,34.152875,-118.486056,0,79.7,0,0,Offer E,13129,0,0,0,0,6,0,0.0,289.92,0.0,497.6,0,1,91436
6838,1,0,0,0,13,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Mailed check,99.0,1301.7,1,31,23,24.14,3493,1,Burbank,0,1,DSL,34.188339,-118.30094199999999,0,102.96,0,0,None,18112,1,1,0,1,13,4,299.0,313.82,0.0,1301.7,0,0,91501
6839,0,0,0,0,11,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,100.75,1129.75,1,45,31,48.64,2229,1,Burbank,1,0,Cable,34.177267,-118.31003,0,104.78,0,0,None,11517,0,0,0,1,11,3,350.0,535.04,0.0,1129.75,0,0,91502
6840,1,0,0,1,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.3,19.3,0,37,0,8.66,4136,0,Burbank,0,1,NA,34.213049,-118.317651,0,19.3,1,0,Offer E,25882,0,0,0,0,1,1,0.0,8.66,0.0,19.3,0,0,91504
6841,1,0,0,0,5,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,55.75,266.95,0,27,41,30.92,4545,0,Burbank,0,1,Fiber Optic,34.174215000000004,-118.345928,0,55.75,0,0,Offer E,29245,1,0,0,1,5,1,109.0,154.60000000000005,0.0,266.95,1,0,91505
6842,1,0,0,0,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Mailed check,19.95,257,0,42,0,16.35,5221,0,Burbank,0,1,NA,34.169706,-118.323548,0,19.95,0,0,None,18539,0,0,0,0,13,0,0.0,212.55,0.0,257.0,0,0,91506
6843,0,0,1,0,9,1,1,Fiber optic,1,1,0,0,Month-to-month,0,Bank transfer (automatic),91.75,865.8,1,58,8,22.0,4176,1,North Hollywood,1,0,Cable,34.1692,-118.372498,1,95.42,0,1,Offer E,36625,0,1,1,0,9,5,0.0,198.0,0.0,865.8,0,1,91601
6844,1,0,0,0,29,1,0,Fiber optic,0,1,1,0,Month-to-month,0,Mailed check,89.65,2623.65,0,39,24,12.92,2681,0,North Hollywood,0,1,DSL,34.15136,-118.36478600000001,0,89.65,0,0,None,16996,1,0,0,0,29,0,0.0,374.68,0.0,2623.65,0,1,91602
6845,1,1,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,45.85,45.85,0,71,6,40.38,5715,0,Studio City,0,1,DSL,34.139082,-118.39275,0,45.85,0,0,None,26157,0,0,0,0,1,1,0.0,40.38,0.0,45.85,0,1,91604
6846,0,0,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,79.55,79.55,1,56,11,5.1,5571,1,North Hollywood,1,0,DSL,34.207295,-118.40002199999999,0,82.73200000000001,0,0,Offer E,57146,0,0,0,0,1,2,0.0,5.1,0.0,79.55,0,0,91605
6847,0,0,1,1,18,1,0,DSL,0,0,1,0,Month-to-month,0,Mailed check,55.95,1082.8,0,33,30,18.47,2035,0,North Hollywood,0,0,DSL,34.187599,-118.387125,1,55.95,4,1,None,45358,0,0,1,0,18,1,0.0,332.46,0.0,1082.8,0,1,91606
6848,0,0,1,0,2,1,0,DSL,0,0,1,1,Month-to-month,0,Credit card (automatic),69.0,147.8,0,61,23,27.41,2798,0,Valley Village,1,0,DSL,34.165783000000005,-118.399795,1,69.0,0,1,Offer E,27453,0,0,1,1,2,0,34.0,54.82,0.0,147.8,0,0,91607
6849,1,0,1,1,30,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),83.55,2570.2,0,19,48,10.24,3558,0,Rancho Cucamonga,0,1,DSL,34.132275,-117.611478,1,83.55,1,1,None,39064,1,0,1,1,30,2,0.0,307.2,0.0,2570.2,1,1,91701
6850,1,0,0,1,66,1,1,DSL,1,1,0,0,Two year,0,Bank transfer (automatic),65.7,4378.9,0,37,17,32.12,5058,0,Azusa,0,1,DSL,34.174493,-117.87068000000001,0,65.7,2,0,None,57775,1,0,0,0,66,0,744.0,2119.92,0.0,4378.9,0,0,91702
6851,1,0,1,1,38,1,1,Fiber optic,0,0,1,0,Two year,1,Bank transfer (automatic),94.9,3616.25,0,32,19,25.84,2436,0,Baldwin Park,1,1,DSL,34.098275,-117.967399,1,94.9,2,1,None,76890,1,0,1,0,38,1,0.0,981.92,0.0,3616.25,0,1,91706
6852,1,0,1,1,44,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,61.9,2924.05,0,41,24,37.68,4388,0,Chino Hills,1,1,Cable,33.942895,-117.72564399999999,1,61.9,3,1,None,66754,1,0,1,0,44,1,70.18,1657.92,0.0,2924.05,0,1,91709
6853,0,0,0,0,54,1,1,Fiber optic,0,1,1,1,Month-to-month,0,Electronic check,111.1,6014.85,1,56,18,46.74,5527,1,Chino,1,0,Cable,33.990646000000005,-117.663025,0,115.544,0,0,None,75319,1,4,0,1,54,3,1083.0,2523.96,0.0,6014.85,0,0,91710
6854,1,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.0,32.7,0,46,0,17.03,3922,0,Claremont,0,1,NA,34.127621000000005,-117.717863,0,20.0,0,0,Offer E,34716,0,0,0,0,2,1,0.0,34.06,0.0,32.7,0,0,91711
6855,0,0,0,0,42,1,0,DSL,1,1,0,1,One year,1,Mailed check,67.7,2882.25,0,55,20,39.32,5034,0,Covina,0,0,Fiber Optic,34.097345000000004,-117.90673600000001,0,67.7,0,0,None,33817,1,0,0,1,42,1,576.0,1651.44,0.0,2882.25,0,0,91722
6856,0,0,1,1,58,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),25.15,1509.9,0,56,0,29.5,6444,0,Covina,0,0,NA,34.084747,-117.886844,1,25.15,2,1,None,17554,0,0,1,0,58,1,0.0,1711.0,0.0,1509.9,0,0,91723
6857,1,0,1,1,58,1,0,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,92.85,5305.05,0,38,24,47.69,4879,0,Covina,0,1,DSL,34.081109999999995,-117.853935,1,92.85,1,1,None,25068,0,0,1,1,58,1,1273.0,2766.02,0.0,5305.05,0,0,91724
6858,0,0,1,1,25,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,89.1,2368.4,1,36,28,23.24,4793,1,Rancho Cucamonga,1,0,Fiber Optic,34.100970000000004,-117.57882,1,92.664,0,1,None,51970,0,2,1,1,25,2,663.0,581.0,0.0,2368.4,0,0,91730
6859,0,0,0,0,71,1,1,Fiber optic,1,1,1,1,Two year,0,Mailed check,111.3,7985.9,0,55,19,49.52,5957,0,El Monte,1,0,Fiber Optic,34.079934,-118.046695,0,111.3,0,0,Offer A,30211,1,0,0,1,71,0,1517.0,3515.92,0.0,7985.9,0,0,91731
6860,0,0,0,0,37,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),101.9,3545.35,1,22,65,24.04,4437,1,El Monte,1,0,DSL,34.074492,-118.01462,0,105.976,0,0,None,62660,0,0,0,1,37,1,0.0,889.48,0.0,3545.35,1,1,91732
6861,0,0,1,1,14,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,91.65,1301,1,61,13,9.13,4304,1,South El Monte,0,0,DSL,34.04622,-118.053753,1,95.316,1,1,None,45645,1,1,1,0,14,2,169.0,127.82,0.0,1301.0,0,0,91733
6862,0,1,0,0,4,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,88.85,372.45,1,69,4,12.86,2754,1,Rancho Cucamonga,1,0,Cable,34.245289,-117.642503,0,92.404,0,0,None,23079,0,3,0,0,4,2,15.0,51.44,0.0,372.45,0,0,91737
6863,0,0,1,0,48,1,1,DSL,1,0,0,0,One year,1,Bank transfer (automatic),60.6,2985.25,0,35,13,44.72,4077,0,Rancho Cucamonga,0,0,Fiber Optic,34.133809,-117.523724,1,60.6,0,1,Offer B,12937,1,0,1,0,48,1,0.0,2146.56,0.0,2985.25,0,1,91739
6864,0,1,0,0,3,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,25.3,77.75,1,80,33,0.0,3542,1,Glendora,0,0,Cable,34.119363,-117.85505900000001,0,26.311999999999998,0,0,None,25135,0,2,0,0,3,3,26.0,0.0,0.0,77.75,0,0,91740
6865,0,0,1,0,8,1,0,DSL,1,0,0,1,Two year,0,Mailed check,65.5,564.35,0,23,41,23.68,2985,0,Glendora,0,0,Fiber Optic,34.14649,-117.84981499999999,1,65.5,0,1,Offer E,24973,1,0,1,1,8,1,231.0,189.44,0.0,564.35,1,0,91741
6866,1,0,0,0,1,1,1,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,95.45,95.45,1,56,2,5.59,5962,1,La Puente,0,1,Cable,34.031441,-117.93643600000001,0,99.26799999999999,0,0,None,84965,0,1,0,1,1,2,0.0,5.59,0.0,95.45,0,0,91744
6867,1,0,0,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.95,1311.75,0,32,0,15.32,6212,0,Hacienda Heights,0,1,NA,33.998471,-117.973758,0,19.95,0,0,Offer A,53686,0,0,0,0,67,0,0.0,1026.44,0.0,1311.75,0,0,91745
6868,1,0,0,0,13,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,91.1,1135.7,1,54,29,5.43,5347,1,La Puente,0,1,DSL,34.038983,-117.991372,0,94.744,0,0,Offer D,30802,0,1,0,1,13,4,32.94,70.59,0.0,1135.7,0,1,91746
6869,0,0,1,1,45,1,0,DSL,0,1,0,0,One year,1,Credit card (automatic),54.15,2319.8,1,60,29,42.04,2761,1,Rowland Heights,0,0,Fiber Optic,33.976753,-117.89736699999999,1,56.316,0,1,None,46342,1,0,1,0,45,2,673.0,1891.8,0.0,2319.8,0,0,91748
6870,1,0,0,0,49,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.6,3720.35,0,39,18,23.82,4516,0,La Verne,0,1,Fiber Optic,34.144703,-117.770299,0,74.6,0,0,Offer B,35530,0,0,0,0,49,0,0.0,1167.18,0.0,3720.35,0,1,91750
6871,0,0,1,0,52,1,1,Fiber optic,0,1,1,0,Month-to-month,0,Bank transfer (automatic),94.6,5025.8,0,60,30,29.23,6212,0,Mira Loma,1,0,DSL,33.999992,-117.535395,1,94.6,0,0,Offer B,18980,0,0,0,0,52,0,0.0,1519.96,0.0,5025.8,0,1,91752
6872,0,0,1,0,63,1,0,Fiber optic,1,0,0,0,One year,1,Credit card (automatic),81.15,5224.5,0,20,46,34.51,5294,0,Monterey Park,1,0,Fiber Optic,34.050321999999994,-118.14703700000001,1,81.15,0,7,Offer B,33280,0,0,1,1,63,2,0.0,2174.13,0.0,5224.5,1,1,91754
6873,0,0,1,1,68,1,1,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),89.05,6185.8,0,50,23,47.91,5001,0,Monterey Park,1,0,DSL,34.049172,-118.115022,1,89.05,1,4,Offer A,26933,1,0,1,1,68,1,0.0,3257.88,0.0,6185.8,0,1,91755
6874,0,0,1,0,31,1,0,DSL,0,0,0,0,Month-to-month,1,Mailed check,49.2,1498.55,0,51,15,1.2,2157,0,Mt Baldy,0,0,DSL,34.231318,-117.66203200000001,1,49.2,0,4,None,47,1,0,1,0,31,1,0.0,37.2,0.0,1498.55,0,1,91759
6875,0,0,1,0,64,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.45,1208.6,0,41,0,19.98,5628,0,Ontario,0,0,NA,34.035602000000004,-117.591528,1,19.45,0,8,Offer B,56280,0,0,1,0,64,0,0.0,1278.72,0.0,1208.6,0,0,91761
6876,0,0,1,0,62,1,0,Fiber optic,1,0,1,1,One year,1,Electronic check,104.3,6613.65,0,37,5,44.95,5905,0,Ontario,1,0,DSL,34.057256,-117.667677,1,104.3,0,5,Offer B,54254,1,0,1,1,62,0,331.0,2786.9,0.0,6613.65,0,0,91762
6877,0,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),69.7,69.7,1,64,28,21.52,4620,1,Montclair,0,0,Cable,34.072121,-117.698319,0,72.488,0,0,None,34447,0,0,0,0,1,4,0.0,21.52,0.0,69.7,0,1,91763
6878,0,0,0,0,6,1,0,Fiber optic,0,0,1,1,Month-to-month,1,Electronic check,89.5,573.3,1,58,28,47.92,2898,1,Ontario,0,0,Cable,34.074087,-117.60561799999999,0,93.08,0,0,Offer E,49474,0,1,0,1,6,4,161.0,287.52,0.0,573.3,0,0,91764
6879,0,0,1,0,21,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,86.05,1818.9,0,40,25,14.81,2937,0,Diamond Bar,0,0,DSL,33.992416,-117.807874,1,86.05,0,7,None,46532,1,0,1,0,21,1,45.47,311.01,0.0,1818.9,0,1,91765
6880,0,0,1,1,72,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),25.2,1787.35,0,64,0,39.3,4382,0,Pomona,0,0,NA,34.042286,-117.756106,1,25.2,3,1,Offer A,69974,0,0,1,0,72,0,0.0,2829.6,0.0,1787.35,0,0,91766
6881,0,0,1,1,32,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Electronic check,35.15,1051.05,0,57,14,0.0,3163,0,Pomona,0,0,Fiber Optic,34.083086,-117.737997,1,35.15,1,3,None,46626,0,0,1,0,32,0,0.0,0.0,0.0,1051.05,0,1,91767
6882,0,1,0,0,71,1,1,Fiber optic,1,1,1,0,One year,1,Credit card (automatic),99.65,7181.25,0,68,12,3.91,5448,0,Pomona,0,0,DSL,34.067932,-117.785168,0,99.65,0,0,Offer A,36057,1,0,0,0,71,0,862.0,277.61,0.0,7181.25,0,0,91768
6883,0,0,0,1,34,1,0,Fiber optic,1,1,1,1,Month-to-month,1,Bank transfer (automatic),105.35,3688.6,0,47,21,32.94,5432,0,Rosemead,1,0,DSL,34.065108,-118.08279099999999,0,105.35,3,0,None,61623,0,0,0,1,34,0,775.0,1119.96,0.0,3688.6,0,0,91770
6884,1,0,1,0,3,0,No phone service,DSL,0,0,0,1,Month-to-month,1,Electronic check,35.15,99.75,1,61,14,0.0,2987,1,San Dimas,0,1,Cable,34.102119,-117.815532,1,36.556,0,1,Offer E,33878,0,2,1,1,3,1,14.0,0.0,0.0,99.75,0,0,91773
6885,1,0,0,1,12,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),73.75,871.4,1,27,65,14.96,2010,1,San Gabriel,0,1,DSL,34.114771999999995,-118.089431,0,76.7,1,0,Offer D,23444,0,0,0,1,12,3,566.0,179.52,0.0,871.4,1,0,91775
6886,0,1,0,0,8,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Electronic check,101.35,780.5,1,78,30,43.98,5546,1,San Gabriel,1,0,Cable,34.089927,-118.09564499999999,0,105.404,0,0,None,38041,0,0,0,0,8,4,234.0,351.84,0.0,780.5,0,0,91776
6887,0,0,1,1,35,1,1,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),24.3,821.6,0,38,0,18.86,5998,0,Temple City,0,0,NA,34.101608,-118.055848,1,24.3,3,5,None,32718,0,0,1,0,35,2,0.0,660.1,0.0,821.6,0,0,91780
6888,0,0,1,1,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,80.7,239.45,0,57,17,23.72,2081,0,Upland,0,0,DSL,34.141146,-117.65558300000001,1,80.7,1,5,Offer E,23331,0,0,1,0,3,1,41.0,71.16,0.0,239.45,0,0,91784
6889,1,0,0,0,3,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Mailed check,89.85,244.45,0,24,59,25.1,4096,0,Upland,1,1,Fiber Optic,34.105493,-117.66093400000001,0,89.85,0,0,None,48827,1,0,0,1,3,3,14.42,75.30000000000003,0.0,244.45,1,1,91786
6890,1,0,0,0,53,1,0,DSL,0,0,0,1,One year,1,Electronic check,61.1,3357.9,0,37,24,4.82,5940,0,Walnut,1,1,DSL,34.018353999999995,-117.85491999999999,0,61.1,0,0,Offer B,45118,0,0,0,1,53,2,0.0,255.46,0.0,3357.9,0,1,91789
6891,0,0,1,0,4,0,No phone service,DSL,1,0,0,0,Month-to-month,1,Electronic check,29.05,129.6,0,40,13,0.0,3306,0,West Covina,0,0,Fiber Optic,34.066964,-117.93700700000001,1,29.05,0,2,Offer E,44099,0,0,1,0,4,2,0.0,0.0,0.0,129.6,0,1,91790
6892,0,0,1,1,48,1,0,Fiber optic,1,0,1,1,One year,1,Bank transfer (automatic),99.7,4977.2,0,53,29,36.18,5921,0,West Covina,1,0,Fiber Optic,34.061634000000005,-117.893169,1,99.7,2,2,Offer B,30458,0,0,1,1,48,0,1443.0,1736.64,0.0,4977.2,0,0,91791
6893,0,0,1,1,6,1,0,DSL,1,1,0,0,Month-to-month,0,Credit card (automatic),55.9,365.35,1,55,22,14.51,4914,1,West Covina,0,0,DSL,34.024405,-117.89872199999999,1,58.136,3,1,Offer E,31622,0,1,1,0,6,2,8.04,87.06,0.0,365.35,0,1,91792
6894,1,1,1,0,3,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,105.9,334.65,1,71,2,41.3,2715,1,Alhambra,1,1,Fiber Optic,34.090925,-118.12816399999998,1,110.136,0,1,None,54382,0,0,1,0,3,2,0.0,123.9,0.0,334.65,0,1,91801
6895,1,0,1,1,54,0,No phone service,DSL,0,0,0,1,Two year,0,Credit card (automatic),46.0,2424.05,0,41,19,0.0,4451,0,Alhambra,1,1,Cable,34.074736,-118.145959,1,46.0,1,0,Offer B,30635,1,0,0,1,54,0,46.06,0.0,0.0,2424.05,0,1,91803
6896,0,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,0,Mailed check,43.95,43.95,1,55,10,34.48,3238,1,Alpine,0,0,DSL,32.827184,-116.70372900000001,0,45.70800000000001,0,0,Offer E,16486,0,0,0,0,1,1,0.0,34.48,0.0,43.95,0,0,91901
6897,1,0,0,0,62,1,0,DSL,0,1,1,1,Month-to-month,1,Bank transfer (automatic),80.4,4981.15,0,49,2,48.72,5157,0,Bonita,1,1,Fiber Optic,32.671170000000004,-117.00232,0,80.4,0,0,Offer B,17389,1,0,0,1,62,1,0.0,3020.64,0.0,4981.15,0,1,91902
6898,1,0,1,1,22,1,0,Fiber optic,0,1,1,1,One year,1,Mailed check,100.05,2090.25,0,36,57,9.05,3274,0,Boulevard,1,1,DSL,32.677096999999996,-116.30499099999999,1,100.05,3,10,None,1509,0,0,1,1,22,0,0.0,199.1,0.0,2090.25,0,1,91905
6899,1,0,0,0,1,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),45.1,45.1,1,27,64,11.06,4884,1,Campo,0,1,Cable,32.673483000000004,-116.47286299999999,0,46.903999999999996,0,0,Offer E,3133,0,0,0,1,1,2,0.0,11.06,0.0,45.1,1,1,91906
6900,1,1,0,0,51,1,0,Fiber optic,0,0,1,1,One year,1,Bank transfer (automatic),94.0,4905.75,0,69,21,4.14,6034,0,Chula Vista,1,1,Fiber Optic,32.636792,-117.05498899999999,0,94.0,0,0,None,74025,0,1,0,1,51,2,0.0,211.14,0.0,4905.75,0,1,91910
6901,0,0,0,0,30,1,1,DSL,0,1,1,0,One year,1,Credit card (automatic),68.95,2038.7,0,37,18,22.64,4403,0,Chula Vista,1,0,Cable,32.607964,-117.059459,0,68.95,0,0,Offer C,71126,0,0,0,0,30,0,0.0,679.2,0.0,2038.7,0,1,91911
6902,0,1,1,0,56,1,1,DSL,1,1,0,0,One year,1,Credit card (automatic),68.45,4014,0,75,18,26.82,4368,0,Chula Vista,1,0,Fiber Optic,32.64164,-116.985026,1,68.45,0,1,None,12884,1,0,1,0,56,0,0.0,1501.92,0.0,4014.0,0,1,91913
6903,1,0,1,0,35,1,1,DSL,0,1,1,0,One year,1,Electronic check,69.0,2441.7,0,50,13,45.97,5283,0,Chula Vista,0,1,Fiber Optic,32.688506,-116.93863200000001,1,69.0,0,6,Offer C,2606,1,0,1,0,35,2,0.0,1608.95,0.0,2441.7,0,1,91914
6904,0,1,0,0,64,0,No phone service,DSL,0,1,1,0,Month-to-month,1,Electronic check,43.85,2751,0,77,21,0.0,6055,0,Chula Vista,0,0,Fiber Optic,32.605012,-116.97595,0,43.85,0,0,None,9278,1,0,0,0,64,0,578.0,0.0,0.0,2751.0,0,0,91915
6905,1,0,0,1,30,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,44.5,1307.8,0,61,17,0.0,5833,0,Descanso,0,1,Fiber Optic,32.912664,-116.63538700000001,0,44.5,1,0,Offer C,1587,0,0,0,1,30,1,222.0,0.0,0.0,1307.8,0,0,91916
6906,0,0,1,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Mailed check,18.7,383.65,0,36,0,2.82,2289,0,Dulzura,0,0,NA,32.622999,-116.687855,1,18.7,3,3,Offer C,727,0,0,1,0,25,0,0.0,70.5,0.0,383.65,0,0,91917
6907,0,0,0,0,41,1,0,Fiber optic,0,0,0,0,Month-to-month,0,Bank transfer (automatic),70.25,2868.05,1,25,45,40.78,3407,1,Guatay,0,0,Cable,32.857946000000005,-116.561917,0,73.06,0,0,None,796,0,0,0,1,41,5,1291.0,1671.98,0.0,2868.05,1,0,91931
6908,1,0,0,1,9,1,0,DSL,0,0,1,0,Month-to-month,0,Electronic check,55.35,449.75,1,40,30,41.02,2688,1,Imperial Beach,0,1,DSL,32.579134,-117.119009,0,57.56399999999999,3,0,Offer E,26662,0,4,0,0,9,3,0.0,369.18,0.0,449.75,0,1,91932
6909,0,0,1,0,1,1,0,DSL,1,1,0,0,Month-to-month,1,Mailed check,53.55,53.55,0,21,59,16.06,4504,0,Jacumba,0,0,DSL,32.649786999999996,-116.2237,1,53.55,0,6,Offer E,699,0,0,1,1,1,3,0.0,16.06,0.0,53.55,1,0,91934
6910,1,0,0,1,70,1,1,Fiber optic,1,1,1,1,Two year,1,Electronic check,114.6,7882.5,0,36,17,26.67,5414,0,Jamul,1,1,Fiber Optic,32.695681,-116.79838600000001,0,114.6,2,0,Offer A,8759,1,0,0,1,70,0,0.0,1866.9,0.0,7882.5,0,1,91935
6911,0,0,1,1,57,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),20.1,1087.7,0,32,0,26.67,5506,0,La Mesa,0,0,NA,32.759327,-116.99726000000001,1,20.1,3,9,Offer B,44652,0,0,1,0,57,1,0.0,1520.19,0.0,1087.7,0,0,91941
6912,1,0,0,0,9,1,1,Fiber optic,0,0,1,0,Month-to-month,1,Electronic check,85.5,791.7,0,35,14,11.5,4867,0,La Mesa,0,1,DSL,32.782501,-117.01611000000001,0,85.5,0,0,Offer E,24005,0,0,0,0,9,1,0.0,103.5,0.0,791.7,0,1,91942
6913,0,0,1,1,69,1,1,Fiber optic,0,1,1,1,One year,1,Bank transfer (automatic),108.75,7493.05,0,45,26,46.45,5874,0,Lemon Grove,1,0,Cable,32.733564,-117.03371299999999,1,108.75,1,5,Offer A,24961,1,0,1,1,69,0,1948.0,3205.05,0.0,7493.05,0,0,91945
6914,1,1,1,0,43,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,103.0,4414.3,1,73,29,17.43,2505,1,Mount Laguna,1,1,Cable,32.830852,-116.444601,1,107.12,0,1,Offer B,81,0,1,1,0,43,2,0.0,749.49,0.0,4414.3,0,1,91948
6915,0,0,1,0,72,1,1,Fiber optic,0,0,1,1,Two year,1,Electronic check,97.85,6841.3,0,57,24,2.56,4508,0,National City,1,0,DSL,32.67102,-117.095235,1,97.85,0,7,Offer A,62355,0,0,1,1,72,0,0.0,184.32,0.0,6841.3,0,1,91950
6916,1,0,0,1,44,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),19.55,819.95,0,48,0,14.37,5860,0,Pine Valley,0,1,NA,32.800671,-116.48336299999998,0,19.55,2,0,Offer B,1604,0,0,0,0,44,1,0.0,632.28,0.0,819.95,0,0,91962
6917,0,0,1,0,72,1,1,Fiber optic,1,1,0,0,Two year,1,Bank transfer (automatic),84.05,6052.25,0,24,52,16.15,5515,0,Potrero,0,0,Fiber Optic,32.619465000000005,-116.59360500000001,1,84.05,0,8,Offer A,905,0,0,1,1,72,0,3147.0,1162.8,0.0,6052.25,1,0,91963
6918,0,0,1,0,33,1,0,Fiber optic,1,0,1,1,One year,1,Electronic check,103.75,3361.05,1,47,26,15.66,3824,1,Spring Valley,1,0,Cable,32.726627,-116.99460800000001,1,107.9,0,1,None,56100,1,0,1,1,33,5,874.0,516.78,0.0,3361.05,0,0,91977
6919,1,0,0,0,54,1,1,Fiber optic,0,0,0,1,Month-to-month,0,Credit card (automatic),89.4,4869.5,0,44,15,35.32,5871,0,Spring Valley,1,1,Cable,32.730264,-116.95096299999999,0,89.4,0,0,Offer B,7863,0,0,0,1,54,3,730.0,1907.28,0.0,4869.5,0,0,91978
6920,1,0,0,1,27,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Credit card (automatic),19.7,509.3,0,48,0,32.28,4052,0,Tecate,0,1,NA,32.587557000000004,-116.636816,0,19.7,1,0,Offer C,91,0,0,0,0,27,2,0.0,871.5600000000002,0.0,509.3,0,0,91980
6921,1,0,0,0,54,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Bank transfer (automatic),79.85,4308.25,0,36,3,7.64,5166,0,Bonsall,0,1,DSL,33.290907000000004,-117.202895,0,79.85,0,0,Offer B,3849,0,0,0,0,54,2,0.0,412.56,0.0,4308.25,0,1,92003
6922,1,0,0,0,3,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Credit card (automatic),74.45,221.1,0,41,5,34.8,3956,0,Borrego Springs,0,1,Fiber Optic,33.200369,-116.19231299999998,0,74.45,0,0,None,2863,0,0,0,0,3,0,11.0,104.4,0.0,221.1,0,0,92004
6923,0,0,1,0,53,1,1,DSL,1,1,0,1,One year,0,Bank transfer (automatic),74.1,3833.95,0,41,4,37.14,5136,0,Cardiff By The Sea,1,0,Cable,33.015865999999995,-117.272254,1,74.1,0,3,Offer B,10375,0,0,1,1,53,3,15.34,1968.42,0.0,3833.95,0,1,92007
6924,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.35,69.35,1,57,29,22.03,2843,1,Carlsbad,0,1,DSL,33.148115999999995,-117.30604299999999,0,72.124,0,0,None,35582,0,1,0,0,1,1,0.0,22.03,0.0,69.35,0,0,92008
6925,1,0,1,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Mailed check,18.8,294.95,0,36,0,14.27,3977,0,Carlsbad,0,1,NA,33.098017999999996,-117.25820300000001,1,18.8,0,5,None,43161,0,1,1,0,15,1,0.0,214.05,0.0,294.95,0,0,92009
6926,0,0,0,0,56,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,73.85,4092.85,1,22,76,35.59,5276,1,Del Mar,0,0,Cable,32.948262,-117.25608600000001,0,76.804,0,0,None,13945,0,0,0,1,56,2,0.0,1993.04,0.0,4092.85,1,1,92014
6927,1,0,1,1,5,1,1,DSL,1,1,0,0,Month-to-month,0,Credit card (automatic),64.4,316.9,0,42,15,17.37,3260,0,El Cajon,0,1,Fiber Optic,32.785165,-116.862648,1,64.4,2,7,None,40995,1,0,1,0,5,0,0.0,86.85000000000002,0.0,316.9,0,1,92019
6928,1,0,1,1,48,1,0,DSL,0,1,0,0,One year,1,Credit card (automatic),55.8,2651.2,0,20,85,38.3,3446,0,El Cajon,1,1,Fiber Optic,32.79697,-116.969082,1,55.8,1,1,Offer B,55277,0,0,1,1,48,2,2254.0,1838.4,0.0,2651.2,1,0,92020
6929,0,0,0,1,25,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Credit card (automatic),20.05,471.7,0,41,0,12.87,2192,0,El Cajon,0,0,NA,32.832706,-116.873258,0,20.05,3,0,Offer C,61872,0,1,0,0,25,1,0.0,321.75,0.0,471.7,0,0,92021
6930,0,0,1,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.15,216.75,1,33,32,15.02,2270,1,Encinitas,0,0,DSL,33.054579,-117.25665,1,78.156,0,1,None,47126,0,0,1,0,3,4,69.0,45.06,0.0,216.75,0,0,92024
6931,1,0,0,0,58,1,0,Fiber optic,1,1,1,1,One year,0,Bank transfer (automatic),99.15,5720.95,0,54,14,32.67,6409,0,Escondido,0,1,DSL,33.081478000000004,-117.03381399999999,0,99.15,0,0,Offer B,49281,0,0,0,1,58,2,801.0,1894.86,0.0,5720.95,0,0,92025
6932,1,0,0,0,10,1,0,DSL,0,0,0,1,Month-to-month,1,Bank transfer (automatic),56.75,503.25,0,23,73,30.3,2037,0,Escondido,0,1,Fiber Optic,33.21846,-117.11691599999999,0,56.75,0,0,None,43436,0,0,0,1,10,1,0.0,303.0,0.0,503.25,1,1,92026
6933,1,0,0,0,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,69.6,69.6,1,27,64,46.21,2072,1,Escondido,0,1,Fiber Optic,33.141265000000004,-116.967221,0,72.384,0,0,None,48690,0,1,0,1,1,1,0.0,46.21,0.0,69.6,1,0,92027
6934,1,0,1,0,71,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),104.15,7365.3,0,27,85,3.86,5973,0,Fallbrook,0,1,DSL,33.362575,-117.299644,1,104.15,0,1,Offer A,42239,1,0,1,1,71,0,6261.0,274.06,0.0,7365.3,1,0,92028
6935,0,0,1,1,65,1,1,Fiber optic,0,1,1,1,Two year,1,Credit card (automatic),110.8,7245.9,0,33,19,45.21,6332,0,Escondido,1,0,Cable,33.079834000000005,-117.134275,1,110.8,2,1,Offer B,17944,1,0,1,1,65,2,0.0,2938.65,0.0,7245.9,0,1,92029
6936,1,0,1,1,5,1,1,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,80.15,385,1,57,21,11.54,5124,1,Julian,0,1,Fiber Optic,32.980678000000005,-116.262854,1,83.35600000000002,1,1,None,3577,0,3,1,0,5,2,81.0,57.7,0.0,385.0,0,0,92036
6937,0,0,0,0,28,0,No phone service,DSL,0,0,0,0,Month-to-month,1,Mailed check,35.75,961.4,0,62,2,0.0,2431,0,La Jolla,1,0,DSL,32.853743,-117.25034,0,35.75,0,0,Offer C,42617,1,0,0,0,28,0,0.0,0.0,0.0,961.4,0,1,92037
6938,0,0,1,1,67,1,1,DSL,0,0,0,1,Two year,1,Bank transfer (automatic),69.9,4615.9,0,46,24,14.83,6079,0,Lakeside,1,0,Fiber Optic,32.909873,-116.906774,1,69.9,1,1,Offer A,42277,1,0,1,1,67,1,0.0,993.61,0.0,4615.9,0,1,92040
6939,1,0,0,0,35,1,0,Fiber optic,1,0,0,1,One year,1,Electronic check,89.2,3251.3,0,60,26,49.61,4446,0,Oceanside,0,1,DSL,33.351059,-117.420557,0,89.2,0,0,Offer C,98239,1,0,0,1,35,2,84.53,1736.35,0.0,3251.3,0,1,92054
6940,0,0,1,1,72,0,No phone service,DSL,1,1,0,1,Two year,0,Credit card (automatic),55.65,3880.05,0,28,59,0.0,5192,0,Oceanside,1,0,DSL,33.194742,-117.29032,1,55.65,3,1,Offer A,52895,1,0,1,1,72,2,2289.0,0.0,0.0,3880.05,1,0,92056
6941,0,0,1,1,61,0,No phone service,DSL,1,1,0,1,One year,1,Bank transfer (automatic),50.7,3088.75,0,25,59,0.0,5024,0,Oceanside,0,0,Fiber Optic,33.254497,-117.28587900000001,1,50.7,1,1,Offer B,46893,1,0,1,1,61,1,182.24,0.0,0.0,3088.75,1,1,92057
6942,1,1,0,0,68,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),20.0,1396,0,66,0,10.48,6136,0,Pala,0,1,NA,33.384345,-117.07261899999999,0,20.0,0,0,Offer A,1831,0,0,0,0,68,0,0.0,712.64,0.0,1396.0,0,0,92059
6943,0,0,1,1,1,0,No phone service,DSL,1,0,0,0,Month-to-month,0,Bank transfer (automatic),30.5,30.5,1,37,21,0.0,5171,1,Palomar Mountain,0,0,Cable,33.309852,-116.82309099999999,1,31.72,1,1,None,234,0,0,1,0,1,4,0.0,0.0,0.0,30.5,0,0,92060
6944,1,0,0,0,3,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.1,53.05,0,49,0,16.32,4905,0,Pauma Valley,0,1,NA,33.313828,-116.940501,0,19.1,0,0,None,2615,0,0,0,0,3,1,0.0,48.96,0.0,53.05,0,0,92061
6945,1,0,1,1,70,1,1,Fiber optic,0,1,1,1,Two year,0,Bank transfer (automatic),98.3,6859.5,1,34,3,29.59,4794,1,Poway,0,1,Cable,32.984395,-117.01345400000001,1,102.23200000000001,0,1,Offer A,47969,0,2,1,1,70,2,0.0,2071.3,0.0,6859.5,0,1,92064
6946,0,0,0,1,48,0,No phone service,DSL,0,1,0,1,Month-to-month,0,Credit card (automatic),45.55,2108.35,0,26,48,0.0,4106,0,Ramona,1,0,Fiber Optic,33.044540999999995,-116.833922,0,45.55,2,0,Offer B,33104,0,1,0,1,48,4,1012.0,0.0,0.0,2108.35,1,0,92065
6947,1,0,1,1,68,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),101.05,6770.5,0,36,18,34.62,5570,0,Ranchita,0,1,Fiber Optic,33.215251,-116.53633,1,101.05,1,10,Offer A,339,0,0,1,1,68,1,1219.0,2354.16,0.0,6770.5,0,0,92066
6948,0,0,0,0,47,1,0,Fiber optic,1,0,1,1,One year,1,Electronic check,103.7,4730.6,0,32,13,2.45,4543,0,Rancho Santa Fe,1,0,Fiber Optic,33.012751,-117.200617,0,103.7,0,0,Offer B,7615,1,0,0,1,47,0,0.0,115.15,0.0,4730.6,0,1,92067
6949,1,0,1,1,32,0,No phone service,DSL,0,0,0,0,One year,1,Mailed check,36.25,1151.05,0,48,53,0.0,2609,0,San Marcos,1,1,DSL,33.162624,-117.17086299999998,1,36.25,3,2,Offer C,52664,1,0,1,0,32,0,610.0,0.0,0.0,1151.05,0,0,92069
6950,0,0,1,1,5,1,0,DSL,1,0,0,0,Month-to-month,1,Mailed check,49.4,232.55,0,54,52,47.06,5756,0,Santa Ysabel,0,0,DSL,33.174725,-116.743329,1,49.4,3,3,None,1143,0,0,1,0,5,0,12.09,235.3,0.0,232.55,0,1,92070
6951,1,0,0,0,49,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Credit card (automatic),19.9,1022.6,0,19,0,6.26,5240,0,Santee,0,1,NA,32.847336,-116.99760500000001,0,19.9,0,0,Offer B,53510,0,0,0,0,49,2,0.0,306.74,0.0,1022.6,1,0,92071
6952,0,0,0,0,48,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Bank transfer (automatic),107.4,5121.3,1,20,52,5.19,4956,1,Solana Beach,1,0,DSL,33.001813,-117.263628,0,111.696,0,0,None,12173,0,1,0,1,48,2,266.31,249.12,0.0,5121.3,1,1,92075
6953,0,1,0,0,13,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,82.0,1127.2,1,79,28,4.45,3363,1,San Marcos,0,0,Fiber Optic,33.119028,-117.166036,0,85.28,0,0,None,6760,0,2,0,0,13,2,316.0,57.85,0.0,1127.2,0,0,92078
6954,1,0,0,0,15,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,19.8,309.4,0,53,0,16.13,2681,0,Valley Center,0,1,NA,33.252829999999996,-116.986079,0,19.8,0,0,None,14575,0,2,0,0,15,2,0.0,241.95,0.0,309.4,0,0,92082
6955,0,0,0,0,12,1,0,DSL,0,0,0,0,Month-to-month,1,Electronic check,45.05,523.1,0,50,12,31.22,5624,0,Vista,0,0,DSL,33.17494,-117.24276100000002,0,45.05,0,0,None,62036,0,0,0,0,12,2,0.0,374.64,0.0,523.1,0,1,92083
6956,1,1,0,0,67,1,1,DSL,1,1,0,0,Two year,1,Bank transfer (automatic),64.55,4250.1,0,79,11,28.88,4494,0,Vista,0,1,DSL,33.22784,-117.200024,0,64.55,0,0,Offer A,44692,1,0,0,0,67,1,468.0,1934.96,0.0,4250.1,0,0,92084
6957,1,0,0,0,9,1,0,Fiber optic,0,0,1,0,Month-to-month,0,Electronic check,86.25,770.5,0,25,59,46.34,4754,0,Warner Springs,0,1,DSL,33.323705,-116.626907,0,86.25,0,0,None,1205,1,0,0,0,9,1,455.0,417.06000000000006,0.0,770.5,1,0,92086
6958,0,0,1,1,13,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),19.75,246.7,0,45,0,5.58,4314,0,Rancho Santa Fe,0,0,NA,32.993559999999995,-117.207121,1,19.75,1,7,None,1072,0,0,1,0,13,0,0.0,72.54,0.0,246.7,0,0,92091
6959,0,0,0,0,38,1,0,Fiber optic,0,0,1,1,One year,1,Mailed check,89.1,3342,0,63,18,30.09,2675,0,San Diego,0,0,Fiber Optic,32.725229999999996,-117.171346,0,89.1,0,0,Offer C,27505,0,0,0,1,38,1,60.16,1143.42,0.0,3342.0,0,1,92101
6960,0,1,1,0,42,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,95.55,3930.6,0,66,12,22.89,4121,0,San Diego,1,0,Fiber Optic,32.716007,-117.11746200000002,1,95.55,0,3,None,47140,0,0,1,0,42,0,472.0,961.38,0.0,3930.6,0,0,92102
6961,0,0,1,0,24,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.4,1747.85,1,55,32,17.73,2325,1,San Diego,0,0,Cable,32.747484,-117.166877,1,78.41600000000003,0,1,None,30202,0,1,1,0,24,2,559.0,425.52,0.0,1747.85,0,0,92103
6962,0,1,1,0,27,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,101.25,2754.45,1,72,14,45.82,4853,1,San Diego,1,0,DSL,32.741499,-117.12740900000001,1,105.3,0,1,None,47689,0,0,1,0,27,0,386.0,1237.14,0.0,2754.45,0,0,92104
6963,1,0,1,1,9,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),102.6,897.75,0,32,30,23.42,4062,0,San Diego,1,1,Fiber Optic,32.741859000000005,-117.09035300000001,1,102.6,3,8,Offer E,73006,0,1,1,1,9,1,26.93,210.78000000000003,0.0,897.75,0,1,92105
6964,0,0,1,0,49,0,No phone service,DSL,0,1,1,1,One year,1,Credit card (automatic),56.3,2780.6,0,51,21,0.0,5913,0,San Diego,0,0,Cable,32.71346,-117.236378,1,56.3,0,1,Offer B,18525,1,0,1,1,49,2,0.0,0.0,0.0,2780.6,0,1,92106
6965,0,1,1,0,61,1,1,Fiber optic,1,1,0,0,Month-to-month,1,Credit card (automatic),94.2,5895.45,0,77,29,33.75,5274,0,San Diego,1,0,Fiber Optic,32.741852,-117.243453,1,94.2,0,1,None,27959,1,0,1,0,61,2,1710.0,2058.75,0.0,5895.45,0,0,92107
6966,1,0,0,1,50,0,No phone service,DSL,1,1,1,0,One year,1,Bank transfer (automatic),43.05,2208.05,0,40,76,0.0,5409,0,San Diego,0,1,Fiber Optic,32.774046000000006,-117.142454,0,43.05,3,0,Offer B,11650,0,0,0,0,50,0,1678.0,0.0,0.0,2208.05,0,0,92108
6967,1,1,0,0,25,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.5,2196.15,1,69,3,18.46,4849,1,San Diego,0,1,Fiber Optic,32.787836,-117.232376,0,93.08,0,0,None,46086,0,1,0,0,25,3,66.0,461.5,0.0,2196.15,0,0,92109
6968,0,1,0,0,22,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Bank transfer (automatic),74.4,1692.6,1,79,25,5.09,2407,1,San Diego,0,0,DSL,32.76501,-117.19938,0,77.376,0,0,None,24169,0,1,0,0,22,3,423.0,111.98,0.0,1692.6,0,0,92110
6969,1,0,0,0,1,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,0,Mailed check,20.5,20.5,1,22,0,19.85,3731,1,San Diego,0,1,NA,32.805518,-117.16905200000001,0,20.5,0,0,None,46828,0,0,0,0,1,3,0.0,19.85,0.0,20.5,1,0,92111
6970,1,0,0,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.35,265.35,1,52,14,47.82,3622,1,San Diego,0,1,Fiber Optic,32.697098,-117.11658700000001,0,77.324,0,0,None,47431,0,2,0,0,4,3,37.0,191.28,0.0,265.35,0,0,92113
6971,0,1,1,0,18,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),99.75,1836.25,1,68,16,25.27,5857,1,San Diego,0,0,Cable,32.707892,-117.05512,1,103.74,0,1,None,66838,1,0,1,0,18,2,29.38,454.86,0.0,1836.25,0,1,92114
6972,0,1,0,0,56,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,111.95,6418.9,1,77,31,19.46,4060,1,San Diego,1,0,Cable,32.762506,-117.07245,0,116.428,0,0,Offer B,56887,1,0,0,0,56,3,1990.0,1089.76,0.0,6418.9,0,0,92115
6973,0,1,1,0,53,1,0,Fiber optic,0,1,1,0,One year,1,Electronic check,94.0,4871.45,0,77,25,47.64,6355,0,San Diego,1,0,Fiber Optic,32.765299,-117.122565,1,94.0,0,1,None,33083,1,0,1,0,53,2,1218.0,2524.92,0.0,4871.45,0,0,92116
6974,0,0,1,0,51,1,1,Fiber optic,0,0,1,1,One year,1,Electronic check,98.85,4947.55,0,34,23,47.72,6034,0,San Diego,1,0,Fiber Optic,32.825086,-117.199424,1,98.85,0,1,Offer B,51213,0,0,1,1,51,0,0.0,2433.72,0.0,4947.55,0,1,92117
6975,0,0,1,1,24,1,1,DSL,1,1,0,0,Two year,0,Electronic check,64.35,1558.65,0,23,85,46.54,5461,0,Coronado,1,0,Cable,32.68674,-117.18661200000001,1,64.35,3,0,Offer C,24093,0,0,0,0,24,2,0.0,1116.96,0.0,1558.65,1,1,92118
6976,0,0,1,0,62,1,0,DSL,1,1,1,0,Two year,1,Credit card (automatic),72.0,4284.2,0,22,59,6.41,6489,0,San Diego,1,0,Cable,32.802959,-117.02709499999999,1,72.0,0,1,Offer B,21866,0,0,1,0,62,2,252.77,397.42,0.0,4284.2,1,1,92119
6977,1,0,0,0,24,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,49.7,1218.25,0,21,59,3.72,2911,0,San Diego,0,1,Fiber Optic,32.807867,-117.060993,0,49.7,0,0,Offer C,25569,0,0,0,0,24,0,719.0,89.28,0.0,1218.25,1,0,92120
6978,0,0,1,1,70,1,1,DSL,1,1,1,0,Two year,0,Electronic check,80.7,5617.95,0,50,16,4.11,4412,0,San Diego,1,0,Cable,32.898613,-117.202937,1,80.7,2,6,Offer A,4258,1,0,1,0,70,0,0.0,287.7000000000001,0.0,5617.95,0,1,92121
6979,1,0,0,1,1,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Mailed check,24.2,24.2,0,64,17,0.0,4276,0,San Diego,0,1,Fiber Optic,32.85723,-117.209774,0,24.2,2,0,Offer E,34902,0,0,0,0,1,1,0.0,0.0,0.0,24.2,0,1,92122
6980,1,1,0,0,16,0,No phone service,DSL,0,1,1,0,Month-to-month,1,Mailed check,39.0,679.85,1,68,26,0.0,5692,1,San Diego,0,1,DSL,32.808814,-117.134694,0,40.56,0,0,None,25232,0,5,0,0,16,1,0.0,0.0,0.0,679.85,0,1,92123
6981,0,0,0,0,8,1,0,DSL,0,1,1,0,Month-to-month,1,Electronic check,65.45,554.45,0,36,16,37.37,5227,0,San Diego,0,0,Fiber Optic,32.827238,-117.08928700000001,0,65.45,0,0,Offer E,30206,1,0,0,0,8,3,0.0,298.96,0.0,554.45,0,1,92124
6982,0,0,1,1,72,1,0,DSL,1,1,0,1,Two year,1,Electronic check,74.35,5237.4,0,61,53,17.21,4874,0,San Diego,1,0,Fiber Optic,32.886925,-117.152162,1,74.35,3,8,Offer A,74232,1,0,1,1,72,0,0.0,1239.12,0.0,5237.4,0,1,92126
6983,0,0,0,0,23,1,0,Fiber optic,0,1,0,0,Month-to-month,0,Bank transfer (automatic),83.2,2032.3,0,23,76,19.96,2061,0,San Diego,1,0,DSL,33.017518,-117.11845600000001,0,83.2,0,0,None,20046,1,0,0,0,23,1,0.0,459.08,23.79,2032.3,1,1,92127
6984,1,0,0,1,31,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Credit card (automatic),25.0,789.2,0,20,51,0.0,4242,0,San Diego,0,1,Cable,33.000269,-117.072093,0,25.0,3,0,Offer C,42733,0,0,0,0,31,1,402.0,0.0,22.4,789.2,1,0,92128
6985,1,0,1,1,37,0,No phone service,DSL,1,0,0,0,One year,1,Electronic check,40.2,1525.35,0,23,52,0.0,2308,0,San Diego,1,1,Fiber Optic,32.961064,-117.13491699999999,1,40.2,2,7,Offer C,47224,1,1,1,0,37,3,793.0,0.0,0.0,1525.35,1,0,92129
6986,0,0,1,0,30,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Credit card (automatic),94.1,2804.45,1,63,26,7.01,5255,1,San Diego,0,0,Fiber Optic,32.957195,-117.202542,1,97.86399999999999,0,1,None,28201,1,0,1,0,30,5,729.0,210.3,0.0,2804.45,0,0,92130
6987,0,1,0,0,35,1,1,Fiber optic,1,1,1,1,One year,1,Electronic check,108.35,3726.15,0,72,3,10.73,5139,0,San Diego,1,0,DSL,32.89325,-117.08709099999999,0,108.35,0,0,Offer C,29283,0,0,0,1,35,0,0.0,375.55,0.0,3726.15,0,1,92131
6988,0,0,1,1,23,1,1,DSL,0,1,1,0,Month-to-month,1,Credit card (automatic),69.5,1652.1,0,60,21,27.49,2159,0,San Diego,0,0,Fiber Optic,32.677716,-117.04766599999999,1,69.5,1,6,None,36351,1,0,1,0,23,1,34.69,632.27,16.89,1652.1,0,1,92139
6989,0,0,1,1,20,1,1,DSL,1,0,1,1,One year,0,Bank transfer (automatic),76.0,1588.75,0,21,59,15.29,4085,0,San Diego,0,0,DSL,32.578103000000006,-117.012975,1,76.0,3,7,None,68776,0,0,1,1,20,2,0.0,305.7999999999999,7.3,1588.75,1,1,92154
6990,1,0,1,0,36,1,0,Fiber optic,1,0,1,1,Month-to-month,1,Electronic check,93.6,3366.05,0,24,41,41.33,2701,0,San Ysidro,0,1,Fiber Optic,32.555828000000005,-117.04007299999999,1,93.6,0,3,Offer C,28488,0,0,1,1,36,1,1380.0,1487.88,16.56,3366.05,1,0,92173
6991,0,0,0,0,8,1,1,Fiber optic,0,0,1,1,Month-to-month,0,Bank transfer (automatic),95.65,778.1,1,53,13,29.66,5335,1,Indio,0,0,Cable,33.713891,-116.237257,0,99.476,0,0,None,56307,0,1,0,1,8,4,0.0,237.28,0.0,778.1,0,1,92201
6992,1,0,1,1,71,1,1,Fiber optic,0,1,1,1,One year,0,Bank transfer (automatic),100.55,7113.75,0,22,59,28.34,5876,0,Indio,0,1,Cable,33.752938,-116.23005500000001,1,100.55,1,1,Offer A,2743,0,0,1,1,71,0,4197.0,2012.14,16.99,7113.75,1,0,92203
6993,0,1,1,0,50,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,88.05,4367.35,1,79,4,37.12,5813,1,Indian Wells,0,0,Cable,33.537646,-116.29108899999999,1,91.572,0,1,Offer B,3873,0,0,1,0,50,1,175.0,1856.0,0.0,4367.35,0,0,92210
6994,0,0,1,1,43,1,1,NA,No internet service,No internet service,No internet service,No internet service,One year,1,Bank transfer (automatic),24.45,993.15,0,59,0,28.03,5119,0,Palm Desert,0,0,NA,33.762759,-116.324817,1,24.45,1,9,Offer B,19702,0,0,1,0,43,0,0.0,1205.29,41.33,993.15,0,0,92211
6995,1,0,0,1,57,1,1,DSL,1,1,1,1,Two year,0,Mailed check,89.55,5012.35,0,55,20,9.36,4260,0,Banning,1,1,Fiber Optic,33.936298,-116.849577,0,89.55,2,0,Offer B,25859,1,0,0,1,57,0,1002.0,533.52,30.45,5012.35,0,0,92220
6996,0,0,1,1,41,1,0,DSL,0,1,0,1,One year,1,Bank transfer (automatic),66.5,2728.6,1,49,31,32.02,2517,1,Beaumont,0,0,Fiber Optic,33.946982,-116.977672,1,69.16,0,1,None,17721,1,0,1,1,41,2,846.0,1312.8200000000004,0.0,2728.6,0,0,92223
6997,0,0,1,0,27,1,0,Fiber optic,0,1,0,0,Month-to-month,1,Electronic check,76.1,2093.4,0,26,59,39.67,3291,0,Blythe,0,0,Cable,33.674583,-114.71611999999999,1,76.1,0,0,Offer C,24659,0,0,0,0,27,1,0.0,1071.09,30.14,2093.4,1,1,92225
6998,0,0,0,0,13,1,0,Fiber optic,0,0,0,1,Month-to-month,1,Electronic check,80.5,1011.8,0,22,27,44.99,3895,0,Brawley,0,0,Cable,33.03933,-115.19185700000001,0,80.5,0,0,None,23394,0,0,0,1,13,0,27.32,584.87,24.99,1011.8,1,1,92227
6999,1,0,0,0,3,0,No phone service,DSL,1,1,0,0,Month-to-month,1,Mailed check,35.45,106.85,1,29,94,0.0,2095,1,Cabazon,0,1,Cable,33.929812,-116.76058,0,36.868,0,0,None,2355,0,0,0,0,3,4,0.0,0.0,0.0,106.85,1,1,92230
7000,0,0,0,0,67,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Electronic check,20.55,1343.4,0,28,0,23.12,5462,0,Calexico,0,0,NA,32.690653999999995,-115.431225,0,20.55,0,0,None,27804,0,0,0,0,67,1,0.0,1549.04,30.53,1343.4,1,0,92231
7001,1,0,0,0,3,1,0,DSL,0,1,0,0,Month-to-month,1,Mailed check,49.9,130.1,1,63,18,46.57,5585,1,Calipatria,0,1,Fiber Optic,33.143826000000004,-115.49748500000001,0,51.896,0,0,None,7857,0,0,0,0,3,4,23.0,139.71,0.0,130.1,0,0,92233
7002,0,0,1,0,64,1,1,Fiber optic,0,1,1,1,Two year,1,Bank transfer (automatic),105.4,6794.75,0,61,18,49.26,4512,0,Cathedral City,0,0,Fiber Optic,33.829583,-116.474131,1,105.4,0,8,Offer B,43141,1,0,1,1,64,1,1223.0,3152.64,32.24,6794.75,0,0,92234
7003,1,0,0,0,26,0,No phone service,DSL,0,0,0,0,Month-to-month,0,Electronic check,35.75,1022.5,0,25,47,0.0,2734,0,Coachella,1,1,Fiber Optic,33.680031,-116.171678,0,35.75,0,0,Offer C,23170,1,0,0,0,26,3,481.0,0.0,0.0,1022.5,1,0,92236
7004,1,0,0,0,38,1,1,Fiber optic,0,1,0,1,Month-to-month,1,Credit card (automatic),95.1,3691.2,0,47,11,6.71,5393,0,Desert Center,1,1,Fiber Optic,33.889604999999996,-115.25700900000001,0,95.1,0,0,Offer C,964,0,0,0,1,38,0,40.6,254.98,0.0,3691.2,0,1,92239
7005,1,0,1,0,23,1,0,NA,No internet service,No internet service,No internet service,No internet service,One year,0,Credit card (automatic),19.3,486.2,0,60,0,36.14,2111,0,Desert Hot Springs,0,1,NA,33.948558,-116.516976,1,19.3,0,3,None,22796,0,0,1,0,23,0,0.0,831.22,0.0,486.2,0,0,92240
7006,1,0,0,0,40,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Credit card (automatic),104.5,4036.85,1,51,16,37.69,2832,1,Desert Hot Springs,1,1,Fiber Optic,33.832799,-116.250973,0,108.68,0,0,None,5529,0,2,0,1,40,3,0.0,1507.6,0.0,4036.85,0,1,92241
7007,1,1,1,0,72,0,No phone service,DSL,1,1,1,1,Two year,1,Bank transfer (automatic),63.1,4685.55,0,78,26,0.0,4933,0,Earp,1,1,DSL,34.137741999999996,-114.36514,1,63.1,0,8,Offer A,1564,1,0,1,1,72,1,0.0,0.0,0.0,4685.55,0,1,92242
7008,0,1,0,0,3,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),75.05,256.25,1,68,33,23.82,3553,1,El Centro,0,0,Cable,32.770393,-115.60915,0,78.05199999999999,0,0,None,43712,0,2,0,0,3,4,85.0,71.46000000000002,0.0,256.25,0,0,92243
7009,1,0,0,0,23,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,81.0,1917.1,1,47,26,18.7,5701,1,Heber,1,1,Cable,32.730583,-115.50108300000001,0,84.24000000000002,0,0,Offer D,3535,0,0,0,0,23,4,498.0,430.1,0.0,1917.1,0,0,92249
7010,0,1,1,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,74.45,74.45,1,73,12,31.27,2394,1,Fallbrook,0,0,DSL,33.362575,-117.299644,1,77.42800000000003,0,1,None,42239,0,0,1,0,1,1,0.0,31.27,0.0,74.45,0,0,92028
7011,0,0,0,0,4,1,0,DSL,1,1,0,0,Month-to-month,1,Mailed check,60.4,272.15,1,28,65,18.03,5730,1,Imperial,0,0,DSL,32.858595,-115.662709,0,62.816,0,0,None,14546,1,2,0,0,4,3,177.0,72.12,0.0,272.15,1,0,92251
7012,0,0,1,0,62,1,1,DSL,1,1,1,1,Two year,1,Electronic check,84.95,5150.55,0,46,28,4.7,6307,0,Joshua Tree,0,0,DSL,34.167235999999995,-116.28151100000001,1,84.95,0,1,Offer B,8141,1,0,1,1,62,0,144.22,291.4000000000001,4.68,5150.55,0,1,92252
7013,0,0,0,0,40,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Bank transfer (automatic),93.4,3756.4,0,54,22,2.83,3819,0,La Quinta,1,0,Cable,33.695532,-116.310571,0,93.4,0,0,Offer B,23971,0,0,0,0,40,2,0.0,113.2,4.18,3756.4,0,1,92253
7014,1,0,0,0,41,1,1,Fiber optic,0,1,1,0,Month-to-month,1,Electronic check,89.2,3645.75,0,35,16,41.85,3259,0,Mecca,0,1,Fiber Optic,33.543834999999994,-115.99390600000001,0,89.2,0,0,Offer B,8768,0,0,0,0,41,0,583.0,1715.85,2.21,3645.75,0,0,92254
7015,1,1,1,0,34,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Credit card (automatic),85.2,2874.45,0,80,29,29.66,5393,0,Morongo Valley,1,1,Cable,34.097863000000004,-116.59456100000001,1,85.2,0,4,Offer C,3499,0,0,1,0,34,0,834.0,1008.44,0.0,2874.45,0,0,92256
7016,0,0,0,0,1,1,0,DSL,0,1,0,0,Month-to-month,0,Electronic check,49.95,49.95,0,37,27,44.98,5230,0,Niland,0,0,Fiber Optic,33.345825,-115.596574,0,49.95,0,0,None,2753,0,0,0,0,1,1,0.0,44.98,0.0,49.95,0,1,92257
7017,0,0,0,0,51,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Bank transfer (automatic),20.65,1020.75,0,25,0,19.23,4725,0,North Palm Springs,0,0,NA,33.906496000000004,-116.569499,0,20.65,0,0,Offer B,732,0,0,0,0,51,1,0.0,980.73,19.32,1020.75,1,0,92258
7018,1,0,1,1,1,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,70.65,70.65,1,64,29,37.68,3463,1,Ocotillo,0,1,DSL,32.698964000000004,-115.886656,1,73.47600000000001,2,1,None,471,0,2,1,0,1,3,0.0,37.68,0.0,70.65,0,1,92259
7019,0,0,0,0,39,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,0,Mailed check,20.15,826,0,30,0,1.57,2007,0,Palm Desert,0,0,NA,33.694501,-116.41271100000002,0,20.15,0,0,Offer C,29340,0,1,0,0,39,1,0.0,61.23,25.92,826.0,0,0,92260
7020,1,0,1,1,12,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Electronic check,19.2,239,0,39,0,25.33,3101,0,Palm Springs,0,1,NA,33.839989,-116.65921499999999,1,19.2,1,2,None,24924,0,0,1,0,12,0,0.0,303.96,45.46,239.0,0,0,92262
7021,1,0,0,0,12,1,0,DSL,0,0,1,0,One year,1,Electronic check,59.8,727.8,1,44,25,9.6,4581,1,Palm Springs,0,1,DSL,33.745746000000004,-116.514215,0,62.192,0,0,Offer D,18884,1,0,0,0,12,3,0.0,115.2,0.0,727.8,0,1,92264
7022,1,0,0,0,72,1,1,Fiber optic,0,1,1,1,One year,1,Electronic check,104.95,7544.3,0,45,18,33.93,5760,0,Palo Verde,1,1,Fiber Optic,33.3249,-114.758334,0,104.95,0,0,None,291,0,1,0,1,72,2,135.8,2442.96,25.42,7544.3,0,1,92266
7023,0,1,1,0,63,1,1,Fiber optic,0,1,1,1,Month-to-month,1,Electronic check,103.5,6479.4,0,77,2,18.14,5187,0,Parker Dam,1,0,Cable,34.273872,-114.192901,1,103.5,0,2,None,131,0,0,1,1,63,0,130.0,1142.82,0.0,6479.4,0,0,92267
7024,1,0,1,0,44,1,1,Fiber optic,1,0,0,0,Month-to-month,1,Credit card (automatic),84.8,3626.35,0,53,10,21.39,2770,0,Pioneertown,1,1,Cable,34.201108000000005,-116.593456,1,84.8,0,2,Offer B,354,0,0,1,0,44,0,36.26,941.16,43.96,3626.35,0,1,92268
7025,0,0,0,0,18,1,1,Fiber optic,0,0,0,1,Month-to-month,1,Bank transfer (automatic),95.05,1679.4,0,51,12,7.42,4524,0,Rancho Mirage,1,0,Fiber Optic,33.763678000000006,-116.429928,0,95.05,0,0,None,12465,1,0,0,1,18,0,202.0,133.56,38.65,1679.4,0,0,92270
7026,0,0,0,0,9,1,0,DSL,0,0,0,0,Month-to-month,1,Bank transfer (automatic),44.2,403.35,1,40,32,41.92,2029,1,Seeley,0,0,Fiber Optic,32.790282,-115.689559,0,45.968,0,0,None,1632,0,1,0,0,9,5,129.0,377.28,0.0,403.35,0,0,92273
7027,1,0,0,0,13,1,0,DSL,0,1,1,1,Month-to-month,0,Mailed check,73.35,931.55,0,64,21,40.99,4645,0,Thermal,0,1,Cable,33.53604,-116.119222,0,73.35,0,0,None,17018,1,0,0,1,13,0,19.56,532.87,49.02,931.55,0,1,92274
7028,0,0,1,0,68,1,0,DSL,0,1,1,0,Two year,0,Bank transfer (automatic),64.1,4326.25,0,23,53,8.62,5553,0,Salton City,0,0,Cable,33.28156,-115.955541,1,64.1,0,2,None,799,1,0,1,0,68,1,229.29,586.16,19.12,4326.25,1,1,92275
7029,0,1,0,0,6,0,No phone service,DSL,0,0,1,1,Month-to-month,1,Electronic check,44.4,263.05,0,75,24,0.0,4611,0,Thousand Palms,0,0,Fiber Optic,33.849263,-116.382778,0,44.4,0,0,None,6242,0,0,0,1,6,0,0.0,0.0,0.0,263.05,0,1,92276
7030,0,0,0,0,2,1,0,NA,No internet service,No internet service,No internet service,No internet service,Month-to-month,1,Mailed check,20.05,39.25,0,57,0,6.85,5191,0,Escondido,0,0,NA,33.141265000000004,-116.967221,0,20.05,0,0,Offer E,48690,0,0,0,0,2,1,0.0,13.7,0.0,39.25,0,0,92027
7031,1,1,1,0,55,1,1,DSL,1,1,0,0,One year,0,Credit card (automatic),60.0,3316.1,0,67,23,9.08,4212,0,Twentynine Palms,0,1,Fiber Optic,34.457829,-116.13958899999999,1,60.0,0,2,None,14104,0,0,1,0,55,1,763.0,499.4,0.0,3316.1,0,0,92278
7032,1,1,0,0,1,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Electronic check,75.75,75.75,1,79,25,8.35,5571,1,Escondido,0,1,Cable,33.141265000000004,-116.967221,0,78.78,0,0,None,48690,0,0,0,0,1,4,0.0,8.35,0.0,75.75,0,0,92027
7033,1,0,0,0,38,1,0,Fiber optic,0,0,0,0,Month-to-month,1,Credit card (automatic),69.5,2625.25,0,63,2,35.04,4591,0,Westmorland,0,1,Fiber Optic,33.03679,-115.60503,0,69.5,0,0,None,2388,0,0,0,0,38,1,53.0,1331.52,20.19,2625.25,0,0,92281
7034,0,0,0,0,67,1,1,Fiber optic,1,1,1,0,Month-to-month,1,Credit card (automatic),102.95,6886.25,1,28,33,37.5,5620,1,White Water,1,0,Fiber Optic,33.972293,-116.654195,0,107.068,0,0,Offer A,805,0,0,0,0,67,5,2272.0,2512.5,0.0,6886.25,1,0,92282
7035,1,0,0,0,19,1,0,Fiber optic,0,0,1,0,Month-to-month,1,Bank transfer (automatic),78.7,1495.1,0,57,13,29.55,2464,0,Winterhaven,0,1,Fiber Optic,32.852947,-114.850784,0,78.7,0,0,None,3663,0,0,0,0,19,0,194.0,561.45,26.84,1495.1,0,0,92283
7036,0,0,0,0,12,0,No phone service,DSL,0,1,1,1,One year,0,Electronic check,60.65,743.3,0,62,24,0.0,3740,0,Yucca Valley,1,0,Fiber Optic,34.159534,-116.42598400000001,0,60.65,0,0,None,20486,1,0,0,1,12,0,17.84,0.0,40.41,743.3,0,1,92284
7037,0,0,0,0,72,1,0,NA,No internet service,No internet service,No internet service,No internet service,Two year,1,Bank transfer (automatic),21.15,1419.4,0,30,0,22.77,5306,0,Landers,0,0,NA,34.341737,-116.53941599999999,0,21.15,0,0,None,2182,0,0,0,0,72,0,0.0,1639.44,19.31,1419.4,0,0,92285
7038,1,0,1,1,24,1,1,DSL,1,0,1,1,One year,1,Mailed check,84.8,1990.5,0,38,24,36.05,2140,0,Adelanto,1,1,DSL,34.667815000000004,-117.53618300000001,1,84.8,2,1,Offer C,18980,1,0,1,1,24,2,0.0,865.1999999999998,48.23,1990.5,0,1,92301
7039,0,0,1,1,72,1,1,Fiber optic,0,1,1,1,One year,1,Credit card (automatic),103.2,7362.9,0,30,59,29.66,5560,0,Amboy,1,0,Cable,34.559882,-115.63716399999998,1,103.2,2,4,None,42,0,0,1,1,72,2,4344.0,2135.52,45.38,7362.9,0,0,92304
7040,0,0,1,1,11,0,No phone service,DSL,1,0,0,0,Month-to-month,1,Electronic check,29.6,346.45,0,32,17,0.0,2793,0,Angelus Oaks,0,0,DSL,34.1678,-116.86433000000001,1,29.6,2,1,None,301,0,0,1,0,11,0,0.0,0.0,27.24,346.45,0,1,92305
7041,1,1,1,0,4,1,1,Fiber optic,0,0,0,0,Month-to-month,1,Mailed check,74.4,306.6,1,75,9,10.61,5839,1,Fallbrook,0,1,DSL,33.362575,-117.299644,1,77.376,0,0,None,42239,0,2,0,0,4,2,28.0,42.44,0.0,306.6,0,0,92028
7042,1,0,0,0,66,1,0,Fiber optic,1,0,1,1,Two year,1,Bank transfer (automatic),105.65,6844.5,0,44,11,30.96,5097,0,Apple Valley,1,1,Fiber Optic,34.424926,-117.184503,0,105.65,0,0,None,28819,1,2,0,1,66,1,0.0,2043.36,0.0,6844.5,0,1,92308
